

module HPSS(






   );
























endmodule