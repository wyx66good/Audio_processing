module sin(
        input wire [9:0]i,
        output reg [15:0] data
   );
always @(*) begin
case(i)
     0   : data= 1999   ; 
     1   : data= 2022   ; 
     2   : data= 2045   ; 
     3   : data= 2067   ; 
     4   : data= 2089   ; 
     5   : data= 2112   ; 
     6   : data= 2134   ; 
     7   : data= 2156   ; 
     8   : data= 2178   ; 
     9   : data= 2200   ; 
     10  : data=  2222  ; 
     11  : data=  2244  ; 
     12  : data=  2265  ; 
     13  : data=  2287  ; 
     14  : data=  2308  ; 
     15  : data=  2329  ; 
     16  : data=  2351  ; 
     17  : data=  2372  ; 
     18  : data=  2393  ; 
     19  : data=  2414  ; 
     20  : data=  2435  ; 
     21  : data=  2455  ; 
     22  : data=  2476  ; 
     23  : data=  2496  ; 
     24  : data=  2517  ; 
     25  : data=  2537  ; 
     26  : data=  2557  ; 
     27  : data=  2577  ; 
     28  : data=  2597  ; 
     29  : data=  2617  ; 
     30  : data=  2637  ; 
     31  : data=  2657  ; 
     32  : data=  2676  ; 
     33  : data=  2695  ; 
     34  : data=  2715  ; 
     35  : data=  2734  ; 
     36  : data=  2753  ; 
     37  : data=  2772  ; 
     38  : data=  2791  ; 
     39  : data=  2809  ; 
     40  : data=  2828  ; 
     41  : data=  2846  ; 
     42  : data=  2865  ; 
     43  : data=  2883  ; 
     44  : data=  2901  ; 
     45  : data=  2919  ; 
     46  : data=  2937  ; 
     47  : data=  2954  ; 
     48  : data=  2972  ; 
     49  : data=  2990  ; 
     50  : data=  3007  ; 
     51  : data=  3024  ; 
     52  : data=  3041  ; 
     53  : data=  3058  ; 
     54  : data=  3075  ; 
     55  : data=  3092  ; 
     56  : data=  3108  ; 
     57  : data=  3124  ; 
     58  : data=  3141  ; 
     59  : data=  3157  ; 
     60  : data=  3173  ; 
     61  : data=  3189  ; 
     62  : data=  3205  ; 
     63  : data=  3220  ; 
     64  : data=  3236  ; 
     65  : data=  3251  ; 
     66  : data=  3266  ; 
     67  : data=  3281  ; 
     68  : data=  3296  ; 
     69  : data=  3311  ; 
     70  : data=  3325  ; 
     71  : data=  3340  ; 
     72  : data=  3354  ; 
     73  : data=  3368  ; 
     74  : data=  3382  ; 
     75  : data=  3396  ; 
     76  : data=  3410  ; 
     77  : data=  3424  ; 
     78  : data=  3437  ; 
     79  : data=  3450  ; 
     80  : data=  3464  ; 
     81  : data=  3477  ; 
     82  : data=  3489  ; 
     83  : data=  3502  ; 
     84  : data=  3515  ; 
     85  : data=  3527  ; 
     86  : data=  3539  ; 
     87  : data=  3552  ; 
     88  : data=  3564  ; 
     89  : data=  3575  ; 
     90  : data=  3587  ; 
     91  : data=  3598  ; 
     92  : data=  3610  ; 
     93  : data=  3621  ; 
     94  : data=  3632  ; 
     95  : data=  3643  ; 
     96  : data=  3654  ; 
     97  : data=  3664  ; 
     98  : data=  3675  ; 
     99  : data=  3685  ; 
     100 : data=   3695 ; 
     101 : data=   3705 ; 
     102 : data=   3715 ; 
     103 : data=   3724 ; 
     104 : data=   3734 ; 
     105 : data=   3743 ; 
     106 : data=   3752 ; 
     107 : data=   3761 ; 
     108 : data=   3770 ; 
     109 : data=   3779 ; 
     110 : data=   3787 ; 
     111 : data=   3796 ; 
     112 : data=   3804 ; 
     113 : data=   3812 ; 
     114 : data=   3820 ; 
     115 : data=   3827 ; 
     116 : data=   3835 ; 
     117 : data=   3842 ; 
     118 : data=   3849 ; 
     119 : data=   3856 ; 
     120 : data=   3863 ; 
     121 : data=   3870 ; 
     122 : data=   3876 ; 
     123 : data=   3883 ; 
     124 : data=   3889 ; 
     125 : data=   3895 ; 
     126 : data=   3901 ; 
     127 : data=   3907 ; 
     128 : data=   3912 ; 
     129 : data=   3917 ; 
     130 : data=   3923 ; 
     131 : data=   3928 ; 
     132 : data=   3933 ; 
     133 : data=   3937 ; 
     134 : data=   3942 ; 
     135 : data=   3946 ; 
     136 : data=   3950 ; 
     137 : data=   3954 ; 
     138 : data=   3958 ; 
     139 : data=   3962 ; 
     140 : data=   3965 ; 
     141 : data=   3969 ; 
     142 : data=   3972 ; 
     143 : data=   3975 ; 
     144 : data=   3978 ; 
     145 : data=   3980 ; 
     146 : data=   3983 ; 
     147 : data=   3985 ; 
     148 : data=   3987 ; 
     149 : data=   3989 ; 
     150 : data=   3991 ; 
     151 : data=   3993 ; 
     152 : data=   3994 ; 
     153 : data=   3995 ; 
     154 : data=   3996 ; 
     155 : data=   3997 ; 
     156 : data=   3998 ; 
     157 : data=   3999 ; 
     158 : data=   3999 ; 
     159 : data=   3999 ; 
     160 : data=   4000 ; 
     161 : data=   3999 ; 
     162 : data=   3999 ; 
     163 : data=   3999 ; 
     164 : data=   3998 ; 
     165 : data=   3997 ; 
     166 : data=   3996 ; 
     167 : data=   3995 ; 
     168 : data=   3994 ; 
     169 : data=   3993 ; 
     170 : data=   3991 ; 
     171 : data=   3989 ; 
     172 : data=   3987 ; 
     173 : data=   3985 ; 
     174 : data=   3983 ; 
     175 : data=   3980 ; 
     176 : data=   3978 ; 
     177 : data=   3975 ; 
     178 : data=   3972 ; 
     179 : data=   3969 ; 
     180 : data=   3965 ; 
     181 : data=   3962 ; 
     182 : data=   3958 ; 
     183 : data=   3954 ; 
     184 : data=   3950 ; 
     185 : data=   3946 ; 
     186 : data=   3942 ; 
     187 : data=   3937 ; 
     188 : data=   3933 ; 
     189 : data=   3928 ; 
     190 : data=   3923 ; 
     191 : data=   3917 ; 
     192 : data=   3912 ; 
     193 : data=   3907 ; 
     194 : data=   3901 ; 
     195 : data=   3895 ; 
     196 : data=   3889 ; 
     197 : data=   3883 ; 
     198 : data=   3876 ; 
     199 : data=   3870 ; 
     200 : data=   3863 ; 
     201 : data=   3856 ; 
     202 : data=   3849 ; 
     203 : data=   3842 ; 
     204 : data=   3835 ; 
     205 : data=   3827 ; 
     206 : data=   3820 ; 
     207 : data=   3812 ; 
     208 : data=   3804 ; 
     209 : data=   3796 ; 
     210 : data=   3787 ; 
     211 : data=   3779 ; 
     212 : data=   3770 ; 
     213 : data=   3761 ; 
     214 : data=   3752 ; 
     215 : data=   3743 ; 
     216 : data=   3734 ; 
     217 : data=   3724 ; 
     218 : data=   3715 ; 
     219 : data=   3705 ; 
     220 : data=   3695 ; 
     221 : data=   3685 ; 
     222 : data=   3675 ; 
     223 : data=   3664 ; 
     224 : data=   3654 ; 
     225 : data=   3643 ; 
     226 : data=   3632 ; 
     227 : data=   3621 ; 
     228 : data=   3610 ; 
     229 : data=   3598 ; 
     230 : data=   3587 ; 
     231 : data=   3575 ; 
     232 : data=   3564 ; 
     233 : data=   3552 ; 
     234 : data=   3539 ; 
     235 : data=   3527 ; 
     236 : data=   3515 ; 
     237 : data=   3502 ; 
     238 : data=   3489 ; 
     239 : data=   3477 ; 
     240 : data=   3464 ; 
     241 : data=   3450 ; 
     242 : data=   3437 ; 
     243 : data=   3424 ; 
     244 : data=   3410 ; 
     245 : data=   3396 ; 
     246 : data=   3382 ; 
     247 : data=   3368 ; 
     248 : data=   3354 ; 
     249 : data=   3340 ; 
     250 : data=   3325 ; 
     251 : data=   3311 ; 
     252 : data=   3296 ; 
     253 : data=   3281 ; 
     254 : data=   3266 ; 
     255 : data=   3251 ; 
     256 : data=   3236 ; 
     257 : data=   3220 ; 
     258 : data=   3205 ; 
     259 : data=   3189 ; 
     260 : data=   3173 ; 
     261 : data=   3157 ; 
     262 : data=   3141 ; 
     263 : data=   3124 ; 
     264 : data=   3108 ; 
     265 : data=   3092 ; 
     266 : data=   3075 ; 
     267 : data=   3058 ; 
     268 : data=   3041 ; 
     269 : data=   3024 ; 
     270 : data=   3007 ; 
     271 : data=   2990 ; 
     272 : data=   2972 ; 
     273 : data=   2954 ; 
     274 : data=   2937 ; 
     275 : data=   2919 ; 
     276 : data=   2901 ; 
     277 : data=   2883 ; 
     278 : data=   2865 ; 
     279 : data=   2846 ; 
     280 : data=   2828 ; 
     281 : data=   2809 ; 
     282 : data=   2791 ; 
     283 : data=   2772 ; 
     284 : data=   2753 ; 
     285 : data=   2734 ; 
     286 : data=   2715 ; 
     287 : data=   2695 ; 
     288 : data=   2676 ; 
     289 : data=   2657 ; 
     290 : data=   2637 ; 
     291 : data=   2617 ; 
     292 : data=   2597 ; 
     293 : data=   2577 ; 
     294 : data=   2557 ; 
     295 : data=   2537 ; 
     296 : data=   2517 ; 
     297 : data=   2496 ; 
     298 : data=   2476 ; 
     299 : data=   2455 ; 
     300 : data=   2435 ; 
     301 : data=   2414 ; 
     302 : data=   2393 ; 
     303 : data=   2372 ; 
     304 : data=   2351 ; 
     305 : data=   2329 ; 
     306 : data=   2308 ; 
     307 : data=   2287 ; 
     308 : data=   2265 ; 
     309 : data=   2244 ; 
     310 : data=   2222 ; 
     311 : data=   2200 ; 
     312 : data=   2178 ; 
     313 : data=   2156 ; 
     314 : data=   2134 ; 
     315 : data=   2112 ; 
     316 : data=   2089 ; 
     317 : data=   2067 ; 
     318 : data=   2045 ; 
     319 : data=   2022 ; 
     320 : data=   1999 ; 
     321 : data=   1977 ; 
     322 : data=   1954 ; 
     323 : data=   1931 ; 
     324 : data=   1908 ; 
     325 : data=   1885 ; 
     326 : data=   1862 ; 
     327 : data=   1839 ; 
     328 : data=   1815 ; 
     329 : data=   1792 ; 
     330 : data=   1769 ; 
     331 : data=   1745 ; 
     332 : data=   1722 ; 
     333 : data=   1698 ; 
     334 : data=   1674 ; 
     335 : data=   1650 ; 
     336 : data=   1626 ; 
     337 : data=   1602 ; 
     338 : data=   1578 ; 
     339 : data=   1554 ; 
     340 : data=   1530 ; 
     341 : data=   1506 ; 
     342 : data=   1482 ; 
     343 : data=   1457 ; 
     344 : data=   1433 ; 
     345 : data=   1409 ; 
     346 : data=   1384 ; 
     347 : data=   1359 ; 
     348 : data=   1335 ; 
     349 : data=   1310 ; 
     350 : data=   1285 ; 
     351 : data=   1260 ; 
     352 : data=   1236 ; 
     353 : data=   1211 ; 
     354 : data=   1186 ; 
     355 : data=   1161 ; 
     356 : data=   1136 ; 
     357 : data=   1110 ; 
     358 : data=   1085 ; 
     359 : data=   1060 ; 
     360 : data=   1035 ; 
     361 : data=   1009 ; 
     362 : data=   984  ; 
     363 : data=   959  ; 
     364 : data=   933  ; 
     365 : data=   908  ; 
     366 : data=   882  ; 
     367 : data=   857  ; 
     368 : data=   831  ; 
     369 : data=   806  ; 
     370 : data=   780  ; 
     371 : data=   754  ; 
     372 : data=   728  ; 
     373 : data=   703  ; 
     374 : data=   677  ; 
     375 : data=   651  ; 
     376 : data=   625  ; 
     377 : data=   599  ; 
     378 : data=   573  ; 
     379 : data=   548  ; 
     380 : data=   522  ; 
     381 : data=   496  ; 
     382 : data=   470  ; 
     383 : data=   444  ; 
     384 : data=   418  ; 
     385 : data=   392  ; 
     386 : data=   366  ; 
     387 : data=   339  ; 
     388 : data=   313  ; 
     389 : data=   287  ; 
     390 : data=   261  ; 
     391 : data=   235  ; 
     392 : data=   209  ; 
     393 : data=   183  ; 
     394 : data=   157  ; 
     395 : data=   130  ; 
     396 : data=   104  ; 
     397 : data=   78   ; 
     398 : data=   52   ; 
     399 : data=   26   ; 
     400 : data=   0    ; 
     401 : data=   -26  ; 
     402 : data=   -52  ; 
     403 : data=   -78  ; 
     404 : data=   -104 ; 
     405 : data=   -130 ; 
     406 : data=   -157 ; 
     407 : data=   -183 ; 
     408 : data=   -209 ; 
     409 : data=   -235 ; 
     410 : data=   -261 ; 
     411 : data=   -287 ; 
     412 : data=   -313 ; 
     413 : data=   -339 ; 
     414 : data=   -366 ; 
     415 : data=   -392 ; 
     416 : data=   -418 ; 
     417 : data=   -444 ; 
     418 : data=   -470 ; 
     419 : data=   -496 ; 
     420 : data=   -522 ; 
     421 : data=   -548 ; 
     422 : data=   -573 ; 
     423 : data=   -599 ; 
     424 : data=   -625 ; 
     425 : data=   -651 ; 
     426 : data=   -677 ; 
     427 : data=   -703 ; 
     428 : data=   -728 ; 
     429 : data=   -754 ; 
     430 : data=   -780 ; 
     431 : data=   -806 ; 
     432 : data=   -831 ; 
     433 : data=   -857 ; 
     434 : data=   -882 ; 
     435 : data=   -908 ; 
     436 : data=   -933 ; 
     437 : data=   -959 ; 
     438 : data=   -984 ; 
     439 : data=   -1009; 
     440 : data=   -1035; 
     441 : data=   -1060; 
     442 : data=   -1085; 
     443 : data=   -1110; 
     444 : data=   -1136; 
     445 : data=   -1161; 
     446 : data=   -1186; 
     447 : data=   -1211; 
     448 : data=   -1236; 
     449 : data=   -1260; 
     450 : data=   -1285; 
     451 : data=   -1310; 
     452 : data=   -1335; 
     453 : data=   -1359; 
     454 : data=   -1384; 
     455 : data=   -1409; 
     456 : data=   -1433; 
     457 : data=   -1457; 
     458 : data=   -1482; 
     459 : data=   -1506; 
     460 : data=   -1530; 
     461 : data=   -1554; 
     462 : data=   -1578; 
     463 : data=   -1602; 
     464 : data=   -1626; 
     465 : data=   -1650; 
     466 : data=   -1674; 
     467 : data=   -1698; 
     468 : data=   -1722; 
     469 : data=   -1745; 
     470 : data=   -1769; 
     471 : data=   -1792; 
     472 : data=   -1815; 
     473 : data=   -1839; 
     474 : data=   -1862; 
     475 : data=   -1885; 
     476 : data=   -1908; 
     477 : data=   -1931; 
     478 : data=   -1954; 
     479 : data=   -1977; 
     480 : data=   -1999; 
     481 : data=   -2022; 
     482 : data=   -2045; 
     483 : data=   -2067; 
     484 : data=   -2089; 
     485 : data=   -2112; 
     486 : data=   -2134; 
     487 : data=   -2156; 
     488 : data=   -2178; 
     489 : data=   -2200; 
     490 : data=   -2222; 
     491 : data=   -2244; 
     492 : data=   -2265; 
     493 : data=   -2287; 
     494 : data=   -2308; 
     495 : data=   -2329; 
     496 : data=   -2351; 
     497 : data=   -2372; 
     498 : data=   -2393; 
     499 : data=   -2414; 
     500 : data=   -2435; 
     501 : data=   -2455; 
     502 : data=   -2476; 
     503 : data=   -2496; 
     504 : data=   -2517; 
     505 : data=   -2537; 
     506 : data=   -2557; 
     507 : data=   -2577; 
     508 : data=   -2597; 
     509 : data=   -2617; 
     510 : data=   -2637; 
     511 : data=   -2657; 
     512 : data=   -2676; 
     513 : data=   -2695; 
     514 : data=   -2715; 
     515 : data=   -2734; 
     516 : data=   -2753; 
     517 : data=   -2772; 
     518 : data=   -2791; 
     519 : data=   -2809; 
     520 : data=   -2828; 
     521 : data=   -2846; 
     522 : data=   -2865; 
     523 : data=   -2883; 
     524 : data=   -2901; 
     525 : data=   -2919; 
     526 : data=   -2937; 
     527 : data=   -2954; 
     528 : data=   -2972; 
     529 : data=   -2990; 
     530 : data=   -3007; 
     531 : data=   -3024; 
     532 : data=   -3041; 
     533 : data=   -3058; 
     534 : data=   -3075; 
     535 : data=   -3092; 
     536 : data=   -3108; 
     537 : data=   -3124; 
     538 : data=   -3141; 
     539 : data=   -3157; 
     540 : data=   -3173; 
     541 : data=   -3189; 
     542 : data=   -3205; 
     543 : data=   -3220; 
     544 : data=   -3236; 
     545 : data=   -3251; 
     546 : data=   -3266; 
     547 : data=   -3281; 
     548 : data=   -3296; 
     549 : data=   -3311; 
     550 : data=   -3325; 
     551 : data=   -3340; 
     552 : data=   -3354; 
     553 : data=   -3368; 
     554 : data=   -3382; 
     555 : data=   -3396; 
     556 : data=   -3410; 
     557 : data=   -3424; 
     558 : data=   -3437; 
     559 : data=   -3450; 
     560 : data=   -3464; 
     561 : data=   -3477; 
     562 : data=   -3489; 
     563 : data=   -3502; 
     564 : data=   -3515; 
     565 : data=   -3527; 
     566 : data=   -3539; 
     567 : data=   -3552; 
     568 : data=   -3564; 
     569 : data=   -3575; 
     570 : data=   -3587; 
     571 : data=   -3598; 
     572 : data=   -3610; 
     573 : data=   -3621; 
     574 : data=   -3632; 
     575 : data=   -3643; 
     576 : data=   -3654; 
     577 : data=   -3664; 
     578 : data=   -3675; 
     579 : data=   -3685; 
     580 : data=   -3695; 
     581 : data=   -3705; 
     582 : data=   -3715; 
     583 : data=   -3724; 
     584 : data=   -3734; 
     585 : data=   -3743; 
     586 : data=   -3752; 
     587 : data=   -3761; 
     588 : data=   -3770; 
     589 : data=   -3779; 
     590 : data=   -3787; 
     591 : data=   -3796; 
     592 : data=   -3804; 
     593 : data=   -3812; 
     594 : data=   -3820; 
     595 : data=   -3827; 
     596 : data=   -3835; 
     597 : data=   -3842; 
     598 : data=   -3849; 
     599 : data=   -3856; 
     600 : data=   -3863; 
     601 : data=   -3870; 
     602 : data=   -3876; 
     603 : data=   -3883; 
     604 : data=   -3889; 
     605 : data=   -3895; 
     606 : data=   -3901; 
     607 : data=   -3907; 
     608 : data=   -3912; 
     609 : data=   -3917; 
     610 : data=   -3923; 
     611 : data=   -3928; 
     612 : data=   -3933; 
     613 : data=   -3937; 
     614 : data=   -3942; 
     615 : data=   -3946; 
     616 : data=   -3950; 
     617 : data=   -3954; 
     618 : data=   -3958; 
     619 : data=   -3962; 
     620 : data=   -3965; 
     621 : data=   -3969; 
     622 : data=   -3972; 
     623 : data=   -3975; 
     624 : data=   -3978; 
     625 : data=   -3980; 
     626 : data=   -3983; 
     627 : data=   -3985; 
     628 : data=   -3987; 
     629 : data=   -3989; 
     630 : data=   -3991; 
     631 : data=   -3993; 
     632 : data=   -3994; 
     633 : data=   -3995; 
     634 : data=   -3996; 
     635 : data=   -3997; 
     636 : data=   -3998; 
     637 : data=   -3999; 
     638 : data=   -3999; 
     639 : data=   -3999; 
     640 : data=   -4000; 
     641 : data=   -3999; 
     642 : data=   -3999; 
     643 : data=   -3999; 
     644 : data=   -3998; 
     645 : data=   -3997; 
     646 : data=   -3996; 
     647 : data=   -3995; 
     648 : data=   -3994; 
     649 : data=   -3993; 
     650 : data=   -3991; 
     651 : data=   -3989; 
     652 : data=   -3987; 
     653 : data=   -3985; 
     654 : data=   -3983; 
     655 : data=   -3980; 
     656 : data=   -3978; 
     657 : data=   -3975; 
     658 : data=   -3972; 
     659 : data=   -3969; 
     660 : data=   -3965; 
     661 : data=   -3962; 
     662 : data=   -3958; 
     663 : data=   -3954; 
     664 : data=   -3950; 
     665 : data=   -3946; 
     666 : data=   -3942; 
     667 : data=   -3937; 
     668 : data=   -3933; 
     669 : data=   -3928; 
     670 : data=   -3923; 
     671 : data=   -3917; 
     672 : data=   -3912; 
     673 : data=   -3907; 
     674 : data=   -3901; 
     675 : data=   -3895; 
     676 : data=   -3889; 
     677 : data=   -3883; 
     678 : data=   -3876; 
     679 : data=   -3870; 
     680 : data=   -3863; 
     681 : data=   -3856; 
     682 : data=   -3849; 
     683 : data=   -3842; 
     684 : data=   -3835; 
     685 : data=   -3827; 
     686 : data=   -3820; 
     687 : data=   -3812; 
     688 : data=   -3804; 
     689 : data=   -3796; 
     690 : data=   -3787; 
     691 : data=   -3779; 
     692 : data=   -3770; 
     693 : data=   -3761; 
     694 : data=   -3752; 
     695 : data=   -3743; 
     696 : data=   -3734; 
     697 : data=   -3724; 
     698 : data=   -3715; 
     699 : data=   -3705; 
     700 : data=   -3695; 
     701 : data=   -3685; 
     702 : data=   -3675; 
     703 : data=   -3664; 
     704 : data=   -3654; 
     705 : data=   -3643; 
     706 : data=   -3632; 
     707 : data=   -3621; 
     708 : data=   -3610; 
     709 : data=   -3598; 
     710 : data=   -3587; 
     711 : data=   -3575; 
     712 : data=   -3564; 
     713 : data=   -3552; 
     714 : data=   -3539; 
     715 : data=   -3527; 
     716 : data=   -3515; 
     717 : data=   -3502; 
     718 : data=   -3489; 
     719 : data=   -3477; 
     720 : data=   -3464; 
     721 : data=   -3450; 
     722 : data=   -3437; 
     723 : data=   -3424; 
     724 : data=   -3410; 
     725 : data=   -3396; 
     726 : data=   -3382; 
     727 : data=   -3368; 
     728 : data=   -3354; 
     729 : data=   -3340; 
     730 : data=   -3325; 
     731 : data=   -3311; 
     732 : data=   -3296; 
     733 : data=   -3281; 
     734 : data=   -3266; 
     735 : data=   -3251; 
     736 : data=   -3236; 
     737 : data=   -3220; 
     738 : data=   -3205; 
     739 : data=   -3189; 
     740 : data=   -3173; 
     741 : data=   -3157; 
     742 : data=   -3141; 
     743 : data=   -3124; 
     744 : data=   -3108; 
     745 : data=   -3092; 
     746 : data=   -3075; 
     747 : data=   -3058; 
     748 : data=   -3041; 
     749 : data=   -3024; 
     750 : data=   -3007; 
     751 : data=   -2990; 
     752 : data=   -2972; 
     753 : data=   -2954; 
     754 : data=   -2937; 
     755 : data=   -2919; 
     756 : data=   -2901; 
     757 : data=   -2883; 
     758 : data=   -2865; 
     759 : data=   -2846; 
     760 : data=   -2828; 
     761 : data=   -2809; 
     762 : data=   -2791; 
     763 : data=   -2772; 
     764 : data=   -2753; 
     765 : data=   -2734; 
     766 : data=   -2715; 
     767 : data=   -2695; 
     768 : data=   -2676; 
     769 : data=   -2657; 
     770 : data=   -2637; 
     771 : data=   -2617; 
     772 : data=   -2597; 
     773 : data=   -2577; 
     774 : data=   -2557; 
     775 : data=   -2537; 
     776 : data=   -2517; 
     777 : data=   -2496; 
     778 : data=   -2476; 
     779 : data=   -2455; 
     780 : data=   -2435; 
     781 : data=   -2414; 
     782 : data=   -2393; 
     783 : data=   -2372; 
     784 : data=   -2351; 
     785 : data=   -2329; 
     786 : data=   -2308; 
     787 : data=   -2287; 
     788 : data=   -2265; 
     789 : data=   -2244; 
     790 : data=   -2222; 
     791 : data=   -2200; 
     792 : data=   -2178; 
     793 : data=   -2156; 
     794 : data=   -2134; 
     795 : data=   -2112; 
     796 : data=   -2089; 
     797 : data=   -2067; 
     798 : data=   -2045; 
     799 : data=   -2022; 
     800 : data=   -1999; 
     801 : data=   -1977; 
     802 : data=   -1954; 
     803 : data=   -1931; 
     804 : data=   -1908; 
     805 : data=   -1885; 
     806 : data=   -1862; 
     807 : data=   -1839; 
     808 : data=   -1815; 
     809 : data=   -1792; 
     810 : data=   -1769; 
     811 : data=   -1745; 
     812 : data=   -1722; 
     813 : data=   -1698; 
     814 : data=   -1674; 
     815 : data=   -1650; 
     816 : data=   -1626; 
     817 : data=   -1602; 
     818 : data=   -1578; 
     819 : data=   -1554; 
     820 : data=   -1530; 
     821 : data=   -1506; 
     822 : data=   -1482; 
     823 : data=   -1457; 
     824 : data=   -1433; 
     825 : data=   -1409; 
     826 : data=   -1384; 
     827 : data=   -1359; 
     828 : data=   -1335; 
     829 : data=   -1310; 
     830 : data=   -1285; 
     831 : data=   -1260; 
     832 : data=   -1236; 
     833 : data=   -1211; 
     834 : data=   -1186; 
     835 : data=   -1161; 
     836 : data=   -1136; 
     837 : data=   -1110; 
     838 : data=   -1085; 
     839 : data=   -1060; 
     840 : data=   -1035; 
     841 : data=   -1009; 
     842 : data=   -984 ; 
     843 : data=   -959 ; 
     844 : data=   -933 ; 
     845 : data=   -908 ; 
     846 : data=   -882 ; 
     847 : data=   -857 ; 
     848 : data=   -831 ; 
     849 : data=   -806 ; 
     850 : data=   -780 ; 
     851 : data=   -754 ; 
     852 : data=   -728 ; 
     853 : data=   -703 ; 
     854 : data=   -677 ; 
     855 : data=   -651 ; 
     856 : data=   -625 ; 
     857 : data=   -599 ; 
     858 : data=   -573 ; 
     859 : data=   -548 ; 
     860 : data=   -522 ; 
     861 : data=   -496 ; 
     862 : data=   -470 ; 
     863 : data=   -444 ; 
     864 : data=   -418 ; 
     865 : data=   -392 ; 
     866 : data=   -366 ; 
     867 : data=   -339 ; 
     868 : data=   -313 ; 
     869 : data=   -287 ; 
     870 : data=   -261 ; 
     871 : data=   -235 ; 
     872 : data=   -209 ; 
     873 : data=   -183 ; 
     874 : data=   -157 ; 
     875 : data=   -130 ; 
     876 : data=   -104 ; 
     877 : data=   -78  ; 
     878 : data=   -52  ; 
     879 : data=   -26  ; 
     880 : data=   0    ; 
     881 : data=   26   ; 
     882 : data=   52   ; 
     883 : data=   78   ; 
     884 : data=   104  ; 
     885 : data=   130  ; 
     886 : data=   157  ; 
     887 : data=   183  ; 
     888 : data=   209  ; 
     889 : data=   235  ; 
     890 : data=   261  ; 
     891 : data=   287  ; 
     892 : data=   313  ; 
     893 : data=   339  ; 
     894 : data=   366  ; 
     895 : data=   392  ; 
     896 : data=   418  ; 
     897 : data=   444  ; 
     898 : data=   470  ; 
     899 : data=   496  ; 
     900 : data=   522  ; 
     901 : data=   548  ; 
     902 : data=   573  ; 
     903 : data=   599  ; 
     904 : data=   625  ; 
     905 : data=   651  ; 
     906 : data=   677  ; 
     907 : data=   703  ; 
     908 : data=   728  ; 
     909 : data=   754  ; 
     910 : data=   780  ; 
     911 : data=   806  ; 
     912 : data=   831  ; 
     913 : data=   857  ; 
     914 : data=   882  ; 
     915 : data=   908  ; 
     916 : data=   933  ; 
     917 : data=   959  ; 
     918 : data=   984  ; 
     919 : data=   1009 ; 
     920 : data=   1035 ; 
     921 : data=   1060 ; 
     922 : data=   1085 ; 
     923 : data=   1110 ; 
     924 : data=   1136 ; 
     925 : data=   1161 ; 
     926 : data=   1186 ; 
     927 : data=   1211 ; 
     928 : data=   1236 ; 
     929 : data=   1260 ; 
     930 : data=   1285 ; 
     931 : data=   1310 ; 
     932 : data=   1335 ; 
     933 : data=   1359 ; 
     934 : data=   1384 ; 
     935 : data=   1409 ; 
     936 : data=   1433 ; 
     937 : data=   1457 ; 
     938 : data=   1482 ; 
     939 : data=   1506 ; 
     940 : data=   1530 ; 
     941 : data=   1554 ; 
     942 : data=   1578 ; 
     943 : data=   1602 ; 
     944 : data=   1626 ; 
     945 : data=   1650 ; 
     946 : data=   1674 ; 
     947 : data=   1698 ; 
     948 : data=   1722 ; 
     949 : data=   1745 ; 
     950 : data=   1769 ; 
     951 : data=   1792 ; 
     952 : data=   1815 ; 
     953 : data=   1839 ; 
     954 : data=   1862 ; 
     955 : data=   1885 ; 
     956 : data=   1908 ; 
     957 : data=   1931 ; 
     958 : data=   1954 ; 
     959 : data=   1977 ; 
     960 : data=   2000 ; 
     961 : data=   2022 ; 
     962 : data=   2045 ; 
     963 : data=   2067 ; 
     964 : data=   2089 ; 
     965 : data=   2112 ; 
     966 : data=   2134 ; 
     967 : data=   2156 ; 
     968 : data=   2178 ; 
     969 : data=   2200 ; 
     970 : data=   2222 ; 
     971 : data=   2244 ; 
     972 : data=   2265 ; 
     973 : data=   2287 ; 
     974 : data=   2308 ; 
     975 : data=   2329 ; 
     976 : data=   2351 ; 
     977 : data=   2372 ; 
     978 : data=   2393 ; 
     979 : data=   2414 ; 
     980 : data=   2435 ; 
     981 : data=   2455 ; 
     982 : data=   2476 ; 
     983 : data=   2496 ; 
     984 : data=   2517 ; 
     985 : data=   2537 ; 
     986 : data=   2557 ; 
     987 : data=   2577 ; 
     988 : data=   2597 ; 
     989 : data=   2617 ; 
     990 : data=   2637 ; 
     991 : data=   2657 ; 
     992 : data=   2676 ; 
     993 : data=   2695 ; 
     994 : data=   2715 ; 
     995 : data=   2734 ; 
     996 : data=   2753 ; 
     997 : data=   2772 ; 
     998 : data=   2791 ; 
     999 : data=   2809 ; 
     1000: data=    2828; 
     1001: data=    2846; 
     1002: data=    2865; 
     1003: data=    2883; 
     1004: data=    2901; 
     1005: data=    2919; 
     1006: data=    2937; 
     1007: data=    2954; 
     1008: data=    2972; 
     1009: data=    2990; 
     1010: data=    3007; 
     1011: data=    3024; 
     1012: data=    3041; 
     1013: data=    3058; 
     1014: data=    3075; 
     1015: data=    3092; 
     1016: data=    3108; 
     1017: data=    3124; 
     1018: data=    3141; 
     1019: data=    3157; 
     1020: data=    3173; 
     1021: data=    3189; 
     1022: data=    3205; 
     1023: data=    3220; 
      default:
            data=    'd0;     

endcase

end



endmodule