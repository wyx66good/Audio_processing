module sin(
        input wire [10:0]i,
        output reg [31:0] data
   );
always @(*) begin
case(i)
   0 :   data=   4432    ;
   1 :   data=   4459    ;
   2 :   data=   4047    ;
   3 :   data=   3762    ;
   4 :   data=   3817    ;
   5 :   data=   3723    ;
   6 :   data=   3426    ;
   7 :   data=   3354    ;
   8 :   data=   3403    ;
   9 :   data=   3166    ;
   10 :  data=  2806     ;
   11 :  data=  2661     ;
   12 :  data=  2574     ;
   13 :  data=  2337     ;
   14 :  data=  2102     ;
   15 :  data=  1928     ;
   16 :  data=  1669     ;
   17 :  data=  1467     ;
   18 :  data=  1536     ;
   19 :  data=  1579     ;
   20 :  data=  1275     ;
   21 :  data=  952      ;
   22 :  data=  915      ;
   23 :  data=  823      ;
   24 :  data=  455      ;
   25 :  data=  172      ;
   26 :  data=  72       ;
   27 :  data=  -200     ;
   28 :  data=  -599     ;
   29 :  data=  -789     ;
   30 :  data=  -941     ;
   31 :  data=  -1293    ;
   32 :  data=  -1506    ;
   33 :  data=  -1370    ;
   34 :  data=  -1328    ;
   35 :  data=  -1610    ;
   36 :  data=  -1877    ;
   37 :  data=  -1973    ;
   38 :  data=  -2082    ;
   39 :  data=  -2229    ;
   40 :  data=  -2408    ;
   41 :  data=  -2772    ;
   42 :  data=  -3159    ;
   43 :  data=  -3208    ;
   44 :  data=  -3104    ;
   45 :  data=  -3276    ;
   46 :  data=  -3482    ;
   47 :  data=  -3308    ;
   48 :  data=  -3121    ;
   49 :  data=  -3409    ;
   50 :  data=  -3785    ;
   51 :  data=  -3768    ;
   52 :  data=  -3741    ;
   53 :  data=  -4134    ;
   54 :  data=  -4539    ;
   55 :  data=  -4508    ;
   56 :  data=  -4327    ;
   57 :  data=  -4312    ;
   58 :  data=  -4262    ;
   59 :  data=  -4051    ;
   60 :  data=  -3923    ;
   61 :  data=  -3975    ;
   62 :  data=  -4078    ;
   63 :  data=  -4215    ;
   64 :  data=  -4362    ;
   65 :  data=  -4390    ;
   66 :  data=  -4376    ;
   67 :  data=  -4477    ;
   68 :  data=  -4499    ;
   69 :  data=  -4276    ;
   70 :  data=  -4134    ;
   71 :  data=  -4244    ;
   72 :  data=  -4190    ;
   73 :  data=  -3831    ;
   74 :  data=  -3663    ;
   75 :  data=  -3843    ;
   76 :  data=  -3934    ;
   77 :  data=  -3811    ;
   78 :  data=  -3774    ;
   79 :  data=  -3815    ;
   80 :  data=  -3723    ;
   81 :  data=  -3613    ;
   82 :  data=  -3640    ;
   83 :  data=  -3621    ;
   84 :  data=  -3393    ;
   85 :  data=  -3134    ;
   86 :  data=  -3089    ;
   87 :  data=  -3270    ;
   88 :  data=  -3466    ;
   89 :  data=  -3441    ;
   90 :  data=  -3203    ;
   91 :  data=  -3045    ;
   92 :  data=  -3131    ;
   93 :  data=  -3210    ;
   94 :  data=  -2977    ;
   95 :  data=  -2561    ;
   96 :  data=  -2414    ;
   97 :  data=  -2656    ;
   98 :  data=  -2839    ;
   99 :  data=  -2655    ;
   100 :  data= -2416    ;
   101 :  data= -2452    ;
   102 :  data= -2578    ;
   103 :  data= -2567    ;
   104 :  data= -2476    ;
   105 :  data= -2315    ;
   106 :  data= -2077    ;
   107 :  data= -1981    ;
   108 :  data= -2080    ;
   109 :  data= -2114    ;
   110 :  data= -2045    ;
   111 :  data= -2011    ;
   112 :  data= -1868    ;
   113 :  data= -1601    ;
   114 :  data= -1573    ;
   115 :  data= -1715    ;
   116 :  data= -1522    ;
   117 :  data= -1154    ;
   118 :  data= -1176    ;
   119 :  data= -1407    ;
   120 :  data= -1405    ;
   121 :  data= -1400    ;
   122 :  data= -1619    ;
   123 :  data= -1691    ;
   124 :  data= -1472    ;
   125 :  data= -1296    ;
   126 :  data= -1204    ;
   127 :  data= -986     ;
   128 :  data= -727     ;
   129 :  data= -500     ;
   130 :  data= -108     ;
   131 :  data= 374      ;
   132 :  data= 559      ;
   133 :  data= 408      ;
   134 :  data= 264      ;
   135 :  data= 250      ;
   136 :  data= 168      ;
   137 :  data= -120     ;
   138 :  data= -512     ;
   139 :  data= -725     ;
   140 :  data= -529     ;
   141 :  data= -61      ;
   142 :  data= 290      ;
   143 :  data= 394      ;
   144 :  data= 524      ;
   145 :  data= 830      ;
   146 :  data= 1024     ;
   147 :  data= 856      ;
   148 :  data= 513      ;
   149 :  data= 306      ;
   150 :  data= 230      ;
   151 :  data= 103      ;
   152 :  data= -81      ;
   153 :  data= -157     ;
   154 :  data= -50      ;
   155 :  data= 61       ;
   156 :  data= -4       ;
   157 :  data= -97      ;
   158 :  data= -2       ;
   159 :  data= 117      ;
   160 :  data= 15       ;
   161 :  data= -157     ;
   162 :  data= -228     ;
   163 :  data= -340     ;
   164 :  data= -479     ;
   165 :  data= -434     ;
   166 :  data= -345     ;
   167 :  data= -410     ;
   168 :  data= -366     ;
   169 :  data= -117     ;
   170 :  data= -73      ;
   171 :  data= -239     ;
   172 :  data= -141     ;
   173 :  data= 93       ;
   174 :  data= -15      ;
   175 :  data= -269     ;
   176 :  data= -249     ;
   177 :  data= -158     ;
   178 :  data= -251     ;
   179 :  data= -322     ;
   180 :  data= -252     ;
   181 :  data= -164     ;
   182 :  data= -46      ;
   183 :  data= 104      ;
   184 :  data= 185      ;
   185 :  data= 316      ;
   186 :  data= 662      ;
   187 :  data= 976      ;
   188 :  data= 966      ;
   189 :  data= 842      ;
   190 :  data= 980      ;
   191 :  data= 1353     ;
   192 :  data= 1600     ;
   193 :  data= 1525     ;
   194 :  data= 1369     ;
   195 :  data= 1442     ;
   196 :  data= 1654     ;
   197 :  data= 1726     ;
   198 :  data= 1673     ;
   199 :  data= 1646     ;
   200 :  data= 1683     ;
   201 :  data= 1899     ;
   202 :  data= 2331     ;
   203 :  data= 2645     ;
   204 :  data= 2678     ;
   205 :  data= 2846     ;
   206 :  data= 3315     ;
   207 :  data= 3605     ;
   208 :  data= 3551     ;
   209 :  data= 3546     ;
   210 :  data= 3645     ;
   211 :  data= 3568     ;
   212 :  data= 3472     ;
   213 :  data= 3643     ;
   214 :  data= 3861     ;
   215 :  data= 3894     ;
   216 :  data= 3978     ;
   217 :  data= 4282     ;
   218 :  data= 4576     ;
   219 :  data= 4694     ;
   220 :  data= 4720     ;
   221 :  data= 4680     ;
   222 :  data= 4559     ;
   223 :  data= 4476     ;
   224 :  data= 4527     ;
   225 :  data= 4631     ;
   226 :  data= 4692     ;
   227 :  data= 4765     ;
   228 :  data= 4926     ;
   229 :  data= 5114     ;
   230 :  data= 5191     ;
   231 :  data= 5108     ;
   232 :  data= 4921     ;
   233 :  data= 4738     ;
   234 :  data= 4693     ;
   235 :  data= 4801     ;
   236 :  data= 4831     ;
   237 :  data= 4636     ;
   238 :  data= 4504     ;
   239 :  data= 4697     ;
   240 :  data= 4858     ;
   241 :  data= 4594     ;
   242 :  data= 4235     ;
   243 :  data= 4197     ;
   244 :  data= 4245     ;
   245 :  data= 4138     ;
   246 :  data= 4149     ;
   247 :  data= 4346     ;
   248 :  data= 4346     ;
   249 :  data= 4133     ;
   250 :  data= 4035     ;
   251 :  data= 3988     ;
   252 :  data= 3739     ;
   253 :  data= 3409     ;
   254 :  data= 3133     ;
   255 :  data= 2851     ;
   256 :  data= 2705     ;
   257 :  data= 2789     ;
   258 :  data= 2720     ;
   259 :  data= 2335     ;
   260 :  data= 2114     ;
   261 :  data= 2216     ;
   262 :  data= 2120     ;
   263 :  data= 1680     ;
   264 :  data= 1394     ;
   265 :  data= 1401     ;
   266 :  data= 1325     ;
   267 :  data= 1064     ;
   268 :  data= 874      ;
   269 :  data= 830      ;
   270 :  data= 769      ;
   271 :  data= 563      ;
   272 :  data= 212      ;
   273 :  data= -166     ;
   274 :  data= -386     ;
   275 :  data= -438     ;
   276 :  data= -573     ;
   277 :  data= -955     ;
   278 :  data= -1325    ;
   279 :  data= -1342    ;
   280 :  data= -1180    ;
   281 :  data= -1263    ;
   282 :  data= -1558    ;
   283 :  data= -1740    ;
   284 :  data= -1853    ;
   285 :  data= -2098    ;
   286 :  data= -2331    ;
   287 :  data= -2441    ;
   288 :  data= -2639    ;
   289 :  data= -2906    ;
   290 :  data= -2950    ;
   291 :  data= -2904    ;
   292 :  data= -3111    ;
   293 :  data= -3364    ;
   294 :  data= -3338    ;
   295 :  data= -3334    ;
   296 :  data= -3670    ;
   297 :  data= -4041    ;
   298 :  data= -4143    ;
   299 :  data= -4140    ;
   300 :  data= -4172    ;
   301 :  data= -4147    ;
   302 :  data= -4110    ;
   303 :  data= -4102    ;
   304 :  data= -3995    ;
   305 :  data= -3852    ;
   306 :  data= -3922    ;
   307 :  data= -4064    ;
   308 :  data= -3988    ;
   309 :  data= -3920    ;
   310 :  data= -4165    ;
   311 :  data= -4401    ;
   312 :  data= -4312    ;
   313 :  data= -4206    ;
   314 :  data= -4322    ;
   315 :  data= -4399    ;
   316 :  data= -4329    ;
   317 :  data= -4310    ;
   318 :  data= -4284    ;
   319 :  data= -4108    ;
   320 :  data= -3941    ;
   321 :  data= -3867    ;
   322 :  data= -3742    ;
   323 :  data= -3635    ;
   324 :  data= -3682    ;
   325 :  data= -3707    ;
   326 :  data= -3603    ;
   327 :  data= -3597    ;
   328 :  data= -3715    ;
   329 :  data= -3720    ;
   330 :  data= -3646    ;
   331 :  data= -3652    ;
   332 :  data= -3596    ;
   333 :  data= -3372    ;
   334 :  data= -3199    ;
   335 :  data= -3220    ;
   336 :  data= -3281    ;
   337 :  data= -3239    ;
   338 :  data= -3140    ;
   339 :  data= -3110    ;
   340 :  data= -3154    ;
   341 :  data= -3109    ;
   342 :  data= -2932    ;
   343 :  data= -2827    ;
   344 :  data= -2840    ;
   345 :  data= -2738    ;
   346 :  data= -2489    ;
   347 :  data= -2362    ;
   348 :  data= -2457    ;
   349 :  data= -2628    ;
   350 :  data= -2719    ;
   351 :  data= -2603    ;
   352 :  data= -2320    ;
   353 :  data= -2152    ;
   354 :  data= -2210    ;
   355 :  data= -2255    ;
   356 :  data= -2153    ;
   357 :  data= -2008    ;
   358 :  data= -1864    ;
   359 :  data= -1732    ;
   360 :  data= -1704    ;
   361 :  data= -1744    ;
   362 :  data= -1677    ;
   363 :  data= -1440    ;
   364 :  data= -1154    ;
   365 :  data= -1075    ;
   366 :  data= -1340    ;
   367 :  data= -1623    ;
   368 :  data= -1567    ;
   369 :  data= -1456    ;
   370 :  data= -1630    ;
   371 :  data= -1687    ;
   372 :  data= -1271    ;
   373 :  data= -762     ;
   374 :  data= -424     ;
   375 :  data= -73      ;
   376 :  data= 208      ;
   377 :  data= 314      ;
   378 :  data= 537      ;
   379 :  data= 780      ;
   380 :  data= 507      ;
   381 :  data= -68      ;
   382 :  data= -257     ;
   383 :  data= -157     ;
   384 :  data= -177     ;
   385 :  data= -117     ;
   386 :  data= 166      ;
   387 :  data= 362      ;
   388 :  data= 469      ;
   389 :  data= 732      ;
   390 :  data= 970      ;
   391 :  data= 966      ;
   392 :  data= 904      ;
   393 :  data= 858      ;
   394 :  data= 661      ;
   395 :  data= 380      ;
   396 :  data= 273      ;
   397 :  data= 401      ;
   398 :  data= 618      ;
   399 :  data= 695      ;
   400 :  data= 505      ;
   401 :  data= 231      ;
   402 :  data= 118      ;
   403 :  data= 135      ;
   404 :  data= 148      ;
   405 :  data= 70       ;
   406 :  data= -152     ;
   407 :  data= -334     ;
   408 :  data= -180     ;
   409 :  data= 124      ;
   410 :  data= 153      ;
   411 :  data= 13       ;
   412 :  data= 28       ;
   413 :  data= 34       ;
   414 :  data= -150     ;
   415 :  data= -262     ;
   416 :  data= -180     ;
   417 :  data= -107     ;
   418 :  data= -47      ;
   419 :  data= 76       ;
   420 :  data= 104      ;
   421 :  data= -3       ;
   422 :  data= -35      ;
   423 :  data= 7        ;
   424 :  data= -40      ;
   425 :  data= -122     ;
   426 :  data= -170     ;
   427 :  data= -273     ;
   428 :  data= -358     ;
   429 :  data= -234     ;
   430 :  data= 30       ;
   431 :  data= 245      ;
   432 :  data= 412      ;
   433 :  data= 607      ;
   434 :  data= 828      ;
   435 :  data= 1042     ;
   436 :  data= 1166     ;
   437 :  data= 1152     ;
   438 :  data= 1107     ;
   439 :  data= 1082     ;
   440 :  data= 960      ;
   441 :  data= 825      ;
   442 :  data= 937      ;
   443 :  data= 1210     ;
   444 :  data= 1362     ;
   445 :  data= 1475     ;
   446 :  data= 1716     ;
   447 :  data= 1882     ;
   448 :  data= 1881     ;
   449 :  data= 2016     ;
   450 :  data= 2342     ;
   451 :  data= 2551     ;
   452 :  data= 2636     ;
   453 :  data= 2817     ;
   454 :  data= 3001     ;
   455 :  data= 3034     ;
   456 :  data= 3066     ;
   457 :  data= 3167     ;
   458 :  data= 3195     ;
   459 :  data= 3178     ;
   460 :  data= 3256     ;
   461 :  data= 3405     ;
   462 :  data= 3616     ;
   463 :  data= 3913     ;
   464 :  data= 4066     ;
   465 :  data= 3901     ;
   466 :  data= 3762     ;
   467 :  data= 3979     ;
   468 :  data= 4281     ;
   469 :  data= 4290     ;
   470 :  data= 4124     ;
   471 :  data= 4104     ;
   472 :  data= 4287     ;
   473 :  data= 4514     ;
   474 :  data= 4603     ;
   475 :  data= 4512     ;
   476 :  data= 4421     ;
   477 :  data= 4504     ;
   478 :  data= 4702     ;
   479 :  data= 4852     ;
   480 :  data= 4913     ;
   481 :  data= 4876     ;
   482 :  data= 4694     ;
   483 :  data= 4423     ;
   484 :  data= 4248     ;
   485 :  data= 4224     ;
   486 :  data= 4218     ;
   487 :  data= 4145     ;
   488 :  data= 4064     ;
   489 :  data= 4038     ;
   490 :  data= 4113     ;
   491 :  data= 4327     ;
   492 :  data= 4479     ;
   493 :  data= 4306     ;
   494 :  data= 4000     ;
   495 :  data= 3996     ;
   496 :  data= 4145     ;
   497 :  data= 3962     ;
   498 :  data= 3558     ;
   499 :  data= 3374     ;
   500 :  data= 3330     ;
   501 :  data= 3140     ;
   502 :  data= 2889     ;
   503 :  data= 2677     ;
   504 :  data= 2435     ;
   505 :  data= 2279     ;
   506 :  data= 2330     ;
   507 :  data= 2349     ;
   508 :  data= 2166     ;
   509 :  data= 1971     ;
   510 :  data= 1862     ;
   511 :  data= 1741     ;
   512 :  data= 1640     ;
   513 :  data= 1545     ;
   514 :  data= 1246     ;
   515 :  data= 816      ;
   516 :  data= 633      ;
   517 :  data= 715      ;
   518 :  data= 690      ;
   519 :  data= 498      ;
   520 :  data= 410      ;
   521 :  data= 396      ;
   522 :  data= 153      ;
   523 :  data= -291     ;
   524 :  data= -632     ;
   525 :  data= -888     ;
   526 :  data= -1292    ;
   527 :  data= -1677    ;
   528 :  data= -1740    ;
   529 :  data= -1652    ;
   530 :  data= -1674    ;
   531 :  data= -1671    ;
   532 :  data= -1590    ;
   533 :  data= -1676    ;
   534 :  data= -1881    ;
   535 :  data= -2014    ;
   536 :  data= -2263    ;
   537 :  data= -2706    ;
   538 :  data= -2972    ;
   539 :  data= -2988    ;
   540 :  data= -3092    ;
   541 :  data= -3269    ;
   542 :  data= -3341    ;
   543 :  data= -3469    ;
   544 :  data= -3666    ;
   545 :  data= -3682    ;
   546 :  data= -3685    ;
   547 :  data= -3964    ;
   548 :  data= -4243    ;
   549 :  data= -4237    ;
   550 :  data= -4168    ;
   551 :  data= -4161    ;
   552 :  data= -4047    ;
   553 :  data= -3836    ;
   554 :  data= -3637    ;
   555 :  data= -3515    ;
   556 :  data= -3637    ;
   557 :  data= -3946    ;
   558 :  data= -4069    ;
   559 :  data= -4055    ;
   560 :  data= -4285    ;
   561 :  data= -4604    ;
   562 :  data= -4622    ;
   563 :  data= -4462    ;
   564 :  data= -4312    ;
   565 :  data= -4094    ;
   566 :  data= -3942    ;
   567 :  data= -3986    ;
   568 :  data= -3961    ;
   569 :  data= -3851    ;
   570 :  data= -3936    ;
   571 :  data= -3984    ;
   572 :  data= -3675    ;
   573 :  data= -3447    ;
   574 :  data= -3619    ;
   575 :  data= -3714    ;
   576 :  data= -3483    ;
   577 :  data= -3302    ;
   578 :  data= -3309    ;
   579 :  data= -3378    ;
   580 :  data= -3533    ;
   581 :  data= -3641    ;
   582 :  data= -3519    ;
   583 :  data= -3437    ;
   584 :  data= -3586    ;
   585 :  data= -3591    ;
   586 :  data= -3328    ;
   587 :  data= -3206    ;
   588 :  data= -3240    ;
   589 :  data= -3067    ;
   590 :  data= -2789    ;
   591 :  data= -2727    ;
   592 :  data= -2746    ;
   593 :  data= -2639    ;
   594 :  data= -2543    ;
   595 :  data= -2561    ;
   596 :  data= -2508    ;
   597 :  data= -2305    ;
   598 :  data= -2110    ;
   599 :  data= -2059    ;
   600 :  data= -2104    ;
   601 :  data= -2145    ;
   602 :  data= -2167    ;
   603 :  data= -2158    ;
   604 :  data= -2045    ;
   605 :  data= -1871    ;
   606 :  data= -1809    ;
   607 :  data= -1845    ;
   608 :  data= -1755    ;
   609 :  data= -1511    ;
   610 :  data= -1333    ;
   611 :  data= -1312    ;
   612 :  data= -1356    ;
   613 :  data= -1389    ;
   614 :  data= -1326    ;
   615 :  data= -1113    ;
   616 :  data= -863     ;
   617 :  data= -672     ;
   618 :  data= -429     ;
   619 :  data= -144     ;
   620 :  data= -35      ;
   621 :  data= -31      ;
   622 :  data= 187      ;
   623 :  data= 472      ;
   624 :  data= 351      ;
   625 :  data= -57      ;
   626 :  data= -197     ;
   627 :  data= -29      ;
   628 :  data= 69       ;
   629 :  data= 63       ;
   630 :  data= 184      ;
   631 :  data= 480      ;
   632 :  data= 889      ;
   633 :  data= 1241     ;
   634 :  data= 1256     ;
   635 :  data= 1038     ;
   636 :  data= 1046     ;
   637 :  data= 1196     ;
   638 :  data= 970      ;
   639 :  data= 538      ;
   640 :  data= 501      ;
   641 :  data= 733      ;
   642 :  data= 769      ;
   643 :  data= 721      ;
   644 :  data= 784      ;
   645 :  data= 756      ;
   646 :  data= 622      ;
   647 :  data= 568      ;
   648 :  data= 454      ;
   649 :  data= 230      ;
   650 :  data= 267      ;
   651 :  data= 541      ;
   652 :  data= 567      ;
   653 :  data= 407      ;
   654 :  data= 516      ;
   655 :  data= 744      ;
   656 :  data= 683      ;
   657 :  data= 498      ;
   658 :  data= 467      ;
   659 :  data= 419      ;
   660 :  data= 239      ;
   661 :  data= 183      ;
   662 :  data= 355      ;
   663 :  data= 518      ;
   664 :  data= 535      ;
   665 :  data= 524      ;
   666 :  data= 572      ;
   667 :  data= 578      ;
   668 :  data= 455      ;
   669 :  data= 279      ;
   670 :  data= 186      ;
   671 :  data= 214      ;
   672 :  data= 323      ;
   673 :  data= 495      ;
   674 :  data= 734      ;
   675 :  data= 1021     ;
   676 :  data= 1309     ;
   677 :  data= 1531     ;
   678 :  data= 1616     ;
   679 :  data= 1549     ;
   680 :  data= 1413     ;
   681 :  data= 1348     ;
   682 :  data= 1379     ;
   683 :  data= 1370     ;
   684 :  data= 1308     ;
   685 :  data= 1389     ;
   686 :  data= 1641     ;
   687 :  data= 1807     ;
   688 :  data= 1824     ;
   689 :  data= 1916     ;
   690 :  data= 2098     ;
   691 :  data= 2193     ;
   692 :  data= 2244     ;
   693 :  data= 2340     ;
   694 :  data= 2412     ;
   695 :  data= 2548     ;
   696 :  data= 2885     ;
   697 :  data= 3140     ;
   698 :  data= 3093     ;
   699 :  data= 3114     ;
   700 :  data= 3394     ;
   701 :  data= 3452     ;
   702 :  data= 3178     ;
   703 :  data= 3156     ;
   704 :  data= 3439     ;
   705 :  data= 3469     ;
   706 :  data= 3355     ;
   707 :  data= 3648     ;
   708 :  data= 4072     ;
   709 :  data= 4041     ;
   710 :  data= 3833     ;
   711 :  data= 3907     ;
   712 :  data= 4001     ;
   713 :  data= 3869     ;
   714 :  data= 3835     ;
   715 :  data= 4024     ;
   716 :  data= 4185     ;
   717 :  data= 4345     ;
   718 :  data= 4598     ;
   719 :  data= 4685     ;
   720 :  data= 4552     ;
   721 :  data= 4523     ;
   722 :  data= 4569     ;
   723 :  data= 4389     ;
   724 :  data= 4176     ;
   725 :  data= 4230     ;
   726 :  data= 4349     ;
   727 :  data= 4332     ;
   728 :  data= 4362     ;
   729 :  data= 4448     ;
   730 :  data= 4346     ;
   731 :  data= 4143     ;
   732 :  data= 4123     ;
   733 :  data= 4256     ;
   734 :  data= 4277     ;
   735 :  data= 4096     ;
   736 :  data= 3922     ;
   737 :  data= 3981     ;
   738 :  data= 4118     ;
   739 :  data= 4031     ;
   740 :  data= 3884     ;
   741 :  data= 3941     ;
   742 :  data= 3905     ;
   743 :  data= 3522     ;
   744 :  data= 3200     ;
   745 :  data= 3137     ;
   746 :  data= 2932     ;
   747 :  data= 2546     ;
   748 :  data= 2368     ;
   749 :  data= 2355     ;
   750 :  data= 2316     ;
   751 :  data= 2403     ;
   752 :  data= 2512     ;
   753 :  data= 2280     ;
   754 :  data= 1875     ;
   755 :  data= 1605     ;
   756 :  data= 1262     ;
   757 :  data= 822      ;
   758 :  data= 732      ;
   759 :  data= 970      ;
   760 :  data= 1082     ;
   761 :  data= 1058     ;
   762 :  data= 1069     ;
   763 :  data= 959      ;
   764 :  data= 671      ;
   765 :  data= 306      ;
   766 :  data= -250     ;
   767 :  data= -970     ;
   768 :  data= -1436    ;
   769 :  data= -1496    ;
   770 :  data= -1430    ;
   771 :  data= -1376    ;
   772 :  data= -1306    ;
   773 :  data= -1289    ;
   774 :  data= -1308    ;
   775 :  data= -1297    ;
   776 :  data= -1414    ;
   777 :  data= -1761    ;
   778 :  data= -2106    ;
   779 :  data= -2299    ;
   780 :  data= -2480    ;
   781 :  data= -2720    ;
   782 :  data= -2913    ;
   783 :  data= -3000    ;
   784 :  data= -3038    ;
   785 :  data= -3089    ;
   786 :  data= -3189    ;
   787 :  data= -3334    ;
   788 :  data= -3515    ;
   789 :  data= -3706    ;
   790 :  data= -3846    ;
   791 :  data= -3900    ;
   792 :  data= -3883    ;
   793 :  data= -3800    ;
   794 :  data= -3690    ;
   795 :  data= -3629    ;
   796 :  data= -3572    ;
   797 :  data= -3458    ;
   798 :  data= -3460    ;
   799 :  data= -3743    ;
   800 :  data= -4097    ;
   801 :  data= -4241    ;
   802 :  data= -4195    ;
   803 :  data= -4091    ;
   804 :  data= -4022    ;
   805 :  data= -4003    ;
   806 :  data= -3908    ;
   807 :  data= -3725    ;
   808 :  data= -3731    ;
   809 :  data= -3944    ;
   810 :  data= -4012    ;
   811 :  data= -3970    ;
   812 :  data= -4132    ;
   813 :  data= -4250    ;
   814 :  data= -3980    ;
   815 :  data= -3660    ;
   816 :  data= -3579    ;
   817 :  data= -3439    ;
   818 :  data= -3177    ;
   819 :  data= -3072    ;
   820 :  data= -3049    ;
   821 :  data= -2973    ;
   822 :  data= -3081    ;
   823 :  data= -3341    ;
   824 :  data= -3406    ;
   825 :  data= -3356    ;
   826 :  data= -3432    ;
   827 :  data= -3472    ;
   828 :  data= -3386    ;
   829 :  data= -3344    ;
   830 :  data= -3239    ;
   831 :  data= -2952    ;
   832 :  data= -2807    ;
   833 :  data= -2927    ;
   834 :  data= -2930    ;
   835 :  data= -2695    ;
   836 :  data= -2468    ;
   837 :  data= -2321    ;
   838 :  data= -2247    ;
   839 :  data= -2322    ;
   840 :  data= -2409    ;
   841 :  data= -2351    ;
   842 :  data= -2340    ;
   843 :  data= -2493    ;
   844 :  data= -2611    ;
   845 :  data= -2651    ;
   846 :  data= -2669    ;
   847 :  data= -2456    ;
   848 :  data= -2000    ;
   849 :  data= -1762    ;
   850 :  data= -1889    ;
   851 :  data= -1965    ;
   852 :  data= -1788    ;
   853 :  data= -1619    ;
   854 :  data= -1662    ;
   855 :  data= -1877    ;
   856 :  data= -2082    ;
   857 :  data= -2026    ;
   858 :  data= -1724    ;
   859 :  data= -1523    ;
   860 :  data= -1502    ;
   861 :  data= -1326    ;
   862 :  data= -921     ;
   863 :  data= -598     ;
   864 :  data= -458     ;
   865 :  data= -378     ;
   866 :  data= -369     ;
   867 :  data= -432     ;
   868 :  data= -439     ;
   869 :  data= -440     ;
   870 :  data= -559     ;
   871 :  data= -638     ;
   872 :  data= -539     ;
   873 :  data= -433     ;
   874 :  data= -350     ;
   875 :  data= -107     ;
   876 :  data= 126      ;
   877 :  data= 53       ;
   878 :  data= -24      ;
   879 :  data= 288      ;
   880 :  data= 648      ;
   881 :  data= 621      ;
   882 :  data= 479      ;
   883 :  data= 515      ;
   884 :  data= 465      ;
   885 :  data= 222      ;
   886 :  data= 106      ;
   887 :  data= 153      ;
   888 :  data= 76       ;
   889 :  data= -86      ;
   890 :  data= -95      ;
   891 :  data= 12       ;
   892 :  data= 109      ;
   893 :  data= 218      ;
   894 :  data= 257      ;
   895 :  data= 107      ;
   896 :  data= -39      ;
   897 :  data= 45       ;
   898 :  data= 198      ;
   899 :  data= 223      ;
   900 :  data= 275      ;
   901 :  data= 418      ;
   902 :  data= 404      ;
   903 :  data= 255      ;
   904 :  data= 299      ;
   905 :  data= 424      ;
   906 :  data= 233      ;
   907 :  data= -69      ;
   908 :  data= 6        ;
   909 :  data= 285      ;
   910 :  data= 308      ;
   911 :  data= 206      ;
   912 :  data= 322      ;
   913 :  data= 577      ;
   914 :  data= 747      ;
   915 :  data= 765      ;
   916 :  data= 617      ;
   917 :  data= 454      ;
   918 :  data= 537      ;
   919 :  data= 773      ;
   920 :  data= 859      ;
   921 :  data= 876      ;
   922 :  data= 1077     ;
   923 :  data= 1350     ;
   924 :  data= 1505     ;
   925 :  data= 1632     ;
   926 :  data= 1762     ;
   927 :  data= 1751     ;
   928 :  data= 1618     ;
   929 :  data= 1523     ;
   930 :  data= 1494     ;
   931 :  data= 1518     ;
   932 :  data= 1649     ;
   933 :  data= 1855     ;
   934 :  data= 2026     ;
   935 :  data= 2143     ;
   936 :  data= 2297     ;
   937 :  data= 2501     ;
   938 :  data= 2657     ;
   939 :  data= 2740     ;
   940 :  data= 2846     ;
   941 :  data= 2976     ;
   942 :  data= 3016     ;
   943 :  data= 3041     ;
   944 :  data= 3205     ;
   945 :  data= 3383     ;
   946 :  data= 3420     ;
   947 :  data= 3452     ;
   948 :  data= 3536     ;
   949 :  data= 3524     ;
   950 :  data= 3491     ;
   951 :  data= 3572     ;
   952 :  data= 3587     ;
   953 :  data= 3527     ;
   954 :  data= 3686     ;
   955 :  data= 3885     ;
   956 :  data= 3767     ;
   957 :  data= 3751     ;
   958 :  data= 4226     ;
   959 :  data= 4536     ;
   960 :  data= 4219     ;
   961 :  data= 3972     ;
   962 :  data= 4223     ;
   963 :  data= 4399     ;
   964 :  data= 4228     ;
   965 :  data= 4110     ;
   966 :  data= 4134     ;
   967 :  data= 4128     ;
   968 :  data= 4216     ;
   969 :  data= 4387     ;
   970 :  data= 4328     ;
   971 :  data= 4127     ;
   972 :  data= 4169     ;
   973 :  data= 4332     ;
   974 :  data= 4228     ;
   975 :  data= 3996     ;
   976 :  data= 3989     ;
   977 :  data= 4066     ;
   978 :  data= 3978     ;
   979 :  data= 3918     ;
   980 :  data= 4025     ;
   981 :  data= 3983     ;
   982 :  data= 3729     ;
   983 :  data= 3729     ;
   984 :  data= 3990     ;
   985 :  data= 3898     ;
   986 :  data= 3431     ;
   987 :  data= 3232     ;
   988 :  data= 3341     ;
   989 :  data= 3250     ;
   990 :  data= 2971     ;
   991 :  data= 2811     ;
   992 :  data= 2641     ;
   993 :  data= 2360     ;
   994 :  data= 2232     ;
   995 :  data= 2275     ;
   996 :  data= 2183     ;
   997 :  data= 1949     ;
   998 :  data= 1784     ;
   999 :  data= 1696     ;
   1000 : data=1607      ;
   1001 : data=1516      ;
   1002 : data=1379      ;
   1003 : data=1171      ;
   1004 : data=1009      ;
   1005 : data=965       ;
   1006 : data=905       ;
   1007 : data=653       ;
   1008 : data=299       ;
   1009 : data=131       ;
   1010 : data=89        ;
   1011 : data=-281      ;
   1012 : data=-947      ;
   1013 : data=-1246     ;
   1014 : data=-1053     ;
   1015 : data=-1004     ;
   1016 : data=-1274     ;
   1017 : data=-1419     ;
   1018 : data=-1390     ;
   1019 : data=-1456     ;
   1020 : data=-1529     ;
   1021 : data=-1580     ;
   1022 : data=-1873     ;
   1023 : data=-2274     ;
   1024 : data=-2391     ;
   1025 : data=-2401     ;
   1026 : data=-2633     ;
   1027 : data=-2861     ;
   1028 : data=-2915     ;
   1029 : data=-3083     ;
   1030 : data=-3347     ;
   1031 : data=-3330     ;
   1032 : data=-3201     ;
   1033 : data=-3409     ;
   1034 : data=-3728     ;
   1035 : data=-3697     ;
   1036 : data=-3543     ;
   1037 : data=-3664     ;
   1038 : data=-3870     ;
   1039 : data=-3905     ;
   1040 : data=-3919     ;
   1041 : data=-3973     ;
   1042 : data=-3900     ;
   1043 : data=-3834     ;
   1044 : data=-3995     ;
   1045 : data=-4135     ;
   1046 : data=-4003     ;
   1047 : data=-3897     ;
   1048 : data=-4046     ;
   1049 : data=-4171     ;
   1050 : data=-4108     ;
   1051 : data=-4093     ;
   1052 : data=-4208     ;
   1053 : data=-4311     ;
   1054 : data=-4378     ;
   1055 : data=-4388     ;
   1056 : data=-4240     ;
   1057 : data=-4047     ;
   1058 : data=-4003     ;
   1059 : data=-3970     ;
   1060 : data=-3757     ;
   1061 : data=-3555     ;
   1062 : data=-3587     ;
   1063 : data=-3701     ;
   1064 : data=-3665     ;
   1065 : data=-3549     ;
   1066 : data=-3544     ;
   1067 : data=-3651     ;
   1068 : data=-3684     ;
   1069 : data=-3575     ;
   1070 : data=-3486     ;
   1071 : data=-3574     ;
   1072 : data=-3726     ;
   1073 : data=-3685     ;
   1074 : data=-3416     ;
   1075 : data=-3190     ;
   1076 : data=-3203     ;
   1077 : data=-3225     ;
   1078 : data=-2968     ;
   1079 : data=-2679     ;
   1080 : data=-2762     ;
   1081 : data=-2991     ;
   1082 : data=-2896     ;
   1083 : data=-2619     ;
   1084 : data=-2539     ;
   1085 : data=-2586     ;
   1086 : data=-2596     ;
   1087 : data=-2583     ;
   1088 : data=-2418     ;
   1089 : data=-2091     ;
   1090 : data=-2009     ;
   1091 : data=-2205     ;
   1092 : data=-2113     ;
   1093 : data=-1723     ;
   1094 : data=-1633     ;
   1095 : data=-1783     ;
   1096 : data=-1726     ;
   1097 : data=-1694     ;
   1098 : data=-1925     ;
   1099 : data=-1936     ;
   1100 : data=-1585     ;
   1101 : data=-1425     ;
   1102 : data=-1459     ;
   1103 : data=-1202     ;
   1104 : data=-827      ;
   1105 : data=-710      ;
   1106 : data=-574      ;
   1107 : data=-247      ;
   1108 : data=-122      ;
   1109 : data=-219      ;
   1110 : data=-152      ;
   1111 : data=-29       ;
   1112 : data=-158      ;
   1113 : data=-313      ;
   1114 : data=-236      ;
   1115 : data=-134      ;
   1116 : data=-126      ;
   1117 : data=-21       ;
   1118 : data=228       ;
   1119 : data=472       ;
   1120 : data=649       ;
   1121 : data=760       ;
   1122 : data=791       ;
   1123 : data=760       ;
   1124 : data=709       ;
   1125 : data=673       ;
   1126 : data=671       ;
   1127 : data=657       ;
   1128 : data=651       ;
   1129 : data=711       ;
   1130 : data=690       ;
   1131 : data=489       ;
   1132 : data=437       ;
   1133 : data=681       ;
   1134 : data=717       ;
   1135 : data=375       ;
   1136 : data=270       ;
   1137 : data=529       ;
   1138 : data=531       ;
   1139 : data=277       ;
   1140 : data=308       ;
   1141 : data=490       ;
   1142 : data=460       ;
   1143 : data=471       ;
   1144 : data=631       ;
   1145 : data=607       ;
   1146 : data=532       ;
   1147 : data=694       ;
   1148 : data=717       ;
   1149 : data=421       ;
   1150 : data=373       ;
   1151 : data=672       ;
   1152 : data=753       ;
   1153 : data=642       ;
   1154 : data=736       ;
   1155 : data=794       ;
   1156 : data=543       ;
   1157 : data=332       ;
   1158 : data=354       ;
   1159 : data=350       ;
   1160 : data=324       ;
   1161 : data=485       ;
   1162 : data=727       ;
   1163 : data=906       ;
   1164 : data=1115      ;
   1165 : data=1376      ;
   1166 : data=1561      ;
   1167 : data=1550      ;
   1168 : data=1340      ;
   1169 : data=1173      ;
   1170 : data=1330      ;
   1171 : data=1600      ;
   1172 : data=1542      ;
   1173 : data=1279      ;
   1174 : data=1285      ;
   1175 : data=1614      ;
   1176 : data=1953      ;
   1177 : data=2060      ;
   1178 : data=1940      ;
   1179 : data=1888      ;
   1180 : data=2153      ;
   1181 : data=2470      ;
   1182 : data=2485      ;
   1183 : data=2387      ;
   1184 : data=2463      ;
   1185 : data=2597      ;
   1186 : data=2722      ;
   1187 : data=2933      ;
   1188 : data=3059      ;
   1189 : data=2987      ;
   1190 : data=3018      ;
   1191 : data=3231      ;
   1192 : data=3287      ;
   1193 : data=3171      ;
   1194 : data=3186      ;
   1195 : data=3330      ;
   1196 : data=3449      ;
   1197 : data=3536      ;
   1198 : data=3516      ;
   1199 : data=3400      ;
               
      default:                 
            data=    'd0;     

endcase

end



endmodule





