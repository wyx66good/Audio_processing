//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2022 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
// Functional description: generates twiddle value
// note: There is no need to use this module in the last stage because w(0) is 1

module ipsxe_fft_exp_rom (
    i_clk       ,
    i_clken     ,
    i_rstn      ,
    i_addr      ,
    o_rdata     , // delay 1
    o_blk_exp
);

parameter   FFT_MODE          = 1       ; // 1: FFT; 0: IFFT
parameter   LOG2_FFT_LEN      = 4       ;   
parameter   INPUT_WIDTH       = 16      ;
parameter   SCALE_MODE        = 0       ; // 1: block floating point; 0: unscaled

localparam  UNSCALED_WIDTH    = INPUT_WIDTH + LOG2_FFT_LEN + 1;
localparam  OUTPUT_WIDTH      = SCALE_MODE ? INPUT_WIDTH : UNSCALED_WIDTH;
                               
input                            i_clk        ;
input                            i_clken      ;
input                            i_rstn       ;
input      [LOG2_FFT_LEN-1:0]    i_addr       ;
output reg [OUTPUT_WIDTH*2-1:0]  o_rdata      ;
output     [4:0]                 o_blk_exp    ; 

// ------------------------------------------------------              
reg        [OUTPUT_WIDTH-1:0]    exp_re_rom [2**LOG2_FFT_LEN-1:0];
reg        [OUTPUT_WIDTH-1:0]    exp_im_rom [2**LOG2_FFT_LEN-1:0];
reg        [4:0]    fft_blk_exp[0:0] ;
reg        [4:0]    ifft_blk_exp [0:0];

initial begin
    if (FFT_MODE) begin
        exp_re_rom[0] = 'h7fffeda;
        exp_re_rom[1] = 'h7fffc2a;
        exp_re_rom[2] = 'h7fff8d3;
        exp_re_rom[3] = 'h7fff70e;
        exp_re_rom[4] = 'hc59a;
        exp_re_rom[5] = 'h7ffea50;
        exp_re_rom[6] = 'h7ffea01;
        exp_re_rom[7] = 'h7ffebf8;
        exp_re_rom[8] = 'h129c3;
        exp_re_rom[9] = 'h7ffd069;
        exp_re_rom[10] = 'h7ffd2cc;
        exp_re_rom[11] = 'h7ffd35b;
        exp_re_rom[12] = 'h5e1e;
        exp_re_rom[13] = 'h7ffbc87;
        exp_re_rom[14] = 'h7ffbac7;
        exp_re_rom[15] = 'h7ffb589;
        exp_re_rom[16] = 'h7ffa8d5;
        exp_re_rom[17] = 'h7ffa744;
        exp_re_rom[18] = 'h7ff9ba7;
        exp_re_rom[19] = 'h7ff87bf;
        exp_re_rom[20] = 'h7fe6361;
        exp_re_rom[21] = 'h7ff9ddb;
        exp_re_rom[22] = 'h7ff7b4b;
        exp_re_rom[23] = 'h7ff4d0a;
        exp_re_rom[24] = 'h7fcbc62;
        exp_re_rom[25] = 'h7ffa6df;
        exp_re_rom[26] = 'h7ff5e00;
        exp_re_rom[27] = 'h7ff0c47;
        exp_re_rom[28] = 'h7fb6192;
        exp_re_rom[29] = 'h7ff937f;
        exp_re_rom[30] = 'h7fefcb9;
        exp_re_rom[31] = 'h7fe1282;
        exp_re_rom[32] = 'h7f0d996;
        exp_re_rom[33] = 'h19864;
        exp_re_rom[34] = 'h4b8d;
        exp_re_rom[35] = 'h7ff9bfb;
        exp_re_rom[36] = 'h7fb9006;
        exp_re_rom[37] = 'h4aa2;
        exp_re_rom[38] = 'h7ff8f7d;
        exp_re_rom[39] = 'h7feb4f7;
        exp_re_rom[40] = 'h7f5fbc7;
        exp_re_rom[41] = 'h18588;
        exp_re_rom[42] = 'h4908;
        exp_re_rom[43] = 'h7ff8aa2;
        exp_re_rom[44] = 'h7fb5a64;
        exp_re_rom[45] = 'h7dab;
        exp_re_rom[46] = 'h7ff764e;
        exp_re_rom[47] = 'h7fe1d4a;
        exp_re_rom[48] = 'h7f0f1a0;
        exp_re_rom[49] = 'h3f02c;
        exp_re_rom[50] = 'h1ea4e;
        exp_re_rom[51] = 'h1712c;
        exp_re_rom[52] = 'h39b03;
        exp_re_rom[53] = 'h7ff42ca;
        exp_re_rom[54] = 'h7ff3373;
        exp_re_rom[55] = 'h7fe4956;
        exp_re_rom[56] = 'h7f51527;
        exp_re_rom[57] = 'h34ae2;
        exp_re_rom[58] = 'h176d6;
        exp_re_rom[59] = 'h103c0;
        exp_re_rom[60] = 'h313a5;
        exp_re_rom[61] = 'h7fe26f1;
        exp_re_rom[62] = 'h7fd99eb;
        exp_re_rom[63] = 'h7faf995;
        exp_re_rom[64] = 'h7e2198e;
        exp_re_rom[65] = 'hc0ecf;
        exp_re_rom[66] = 'h668b6;
        exp_re_rom[67] = 'h5ab3a;
        exp_re_rom[68] = 'hc7dd1;
        exp_re_rom[69] = 'h7fefb24;
        exp_re_rom[70] = 'hc038;
        exp_re_rom[71] = 'h135f3;
        exp_re_rom[72] = 'h24da8;
        exp_re_rom[73] = 'h94f0;
        exp_re_rom[74] = 'he7c0;
        exp_re_rom[75] = 'h10f27;
        exp_re_rom[76] = 'h1c1c1;
        exp_re_rom[77] = 'h85d9;
        exp_re_rom[78] = 'hc02a;
        exp_re_rom[79] = 'hd3bd;
        exp_re_rom[80] = 'hf9be;
        exp_re_rom[81] = 'hcc04;
        exp_re_rom[82] = 'he548;
        exp_re_rom[83] = 'h10d8a;
        exp_re_rom[84] = 'h221eb;
        exp_re_rom[85] = 'h7fff4d8;
        exp_re_rom[86] = 'h5602;
        exp_re_rom[87] = 'h5012;
        exp_re_rom[88] = 'h7ff65e4;
        exp_re_rom[89] = 'h17188;
        exp_re_rom[90] = 'h1071c;
        exp_re_rom[91] = 'hcc95;
        exp_re_rom[92] = 'h7ff2af7;
        exp_re_rom[93] = 'h351dc;
        exp_re_rom[94] = 'h3183e;
        exp_re_rom[95] = 'h46e89;
        exp_re_rom[96] = 'he00bb;
        exp_re_rom[97] = 'h7f8dadc;
        exp_re_rom[98] = 'h7fe08b0;
        exp_re_rom[99] = 'h113e;
        exp_re_rom[100] = 'h6f92e;
        exp_re_rom[101] = 'h7f7730c;
        exp_re_rom[102] = 'h7fa8902;
        exp_re_rom[103] = 'h7f989a5;
        exp_re_rom[104] = 'h7ee6560;
        exp_re_rom[105] = 'ha241f;
        exp_re_rom[106] = 'h32ae5;
        exp_re_rom[107] = 'h1693a;
        exp_re_rom[108] = 'h7ff15b7;
        exp_re_rom[109] = 'h33070;
        exp_re_rom[110] = 'h201bd;
        exp_re_rom[111] = 'h21c79;
        exp_re_rom[112] = 'h4f41f;
        exp_re_rom[113] = 'h7fca929;
        exp_re_rom[114] = 'h7feb142;
        exp_re_rom[115] = 'h7fef695;
        exp_re_rom[116] = 'h7ff4db7;
        exp_re_rom[117] = 'h7fd3cd1;
        exp_re_rom[118] = 'h7fc8dd2;
        exp_re_rom[119] = 'h7f9db76;
        exp_re_rom[120] = 'h7eaf4bd;
        exp_re_rom[121] = 'h14a88e;
        exp_re_rom[122] = 'h7d586;
        exp_re_rom[123] = 'h4edce;
        exp_re_rom[124] = 'h1bce4;
        exp_re_rom[125] = 'h86d82;
        exp_re_rom[126] = 'h6bc55;
        exp_re_rom[127] = 'h82798;
        exp_re_rom[128] = 'h12b0c1;
        exp_re_rom[129] = 'h7f0e274;
        exp_re_rom[130] = 'h7fb6c0b;
        exp_re_rom[131] = 'h7fc57cb;
        exp_re_rom[132] = 'h7f6df49;
        exp_re_rom[133] = 'hc755b;
        exp_re_rom[134] = 'h63e03;
        exp_re_rom[135] = 'h6bd9b;
        exp_re_rom[136] = 'he7337;
        exp_re_rom[137] = 'h7f35fc2;
        exp_re_rom[138] = 'h7fd073b;
        exp_re_rom[139] = 'h7fed8d4;
        exp_re_rom[140] = 'h7ffd270;
        exp_re_rom[141] = 'h7ff67ff;
        exp_re_rom[142] = 'h7ffff35;
        exp_re_rom[143] = 'h4c24;
        exp_re_rom[144] = 'hc506;
        exp_re_rom[145] = 'h7ffc051;
        exp_re_rom[146] = 'h4ec0;
        exp_re_rom[147] = 'h838c;
        exp_re_rom[148] = 'he651;
        exp_re_rom[149] = 'h7ffb30f;
        exp_re_rom[150] = 'h21b2;
        exp_re_rom[151] = 'h7fff17d;
        exp_re_rom[152] = 'h7fe69cb;
        exp_re_rom[153] = 'h54af3;
        exp_re_rom[154] = 'h2abce;
        exp_re_rom[155] = 'h28a0c;
        exp_re_rom[156] = 'h348ae;
        exp_re_rom[157] = 'h9aac;
        exp_re_rom[158] = 'h26630;
        exp_re_rom[159] = 'h3cb51;
        exp_re_rom[160] = 'h8d9d1;
        exp_re_rom[161] = 'h7f35924;
        exp_re_rom[162] = 'h7fd57da;
        exp_re_rom[163] = 'h7ff1c34;
        exp_re_rom[164] = 'h8c2d;
        exp_re_rom[165] = 'h7fd35a5;
        exp_re_rom[166] = 'h7ff168b;
        exp_re_rom[167] = 'h7ff3bf3;
        exp_re_rom[168] = 'h7fe05f6;
        exp_re_rom[169] = 'h62bbe;
        exp_re_rom[170] = 'h2d511;
        exp_re_rom[171] = 'h3131f;
        exp_re_rom[172] = 'h55f83;
        exp_re_rom[173] = 'h7fa1216;
        exp_re_rom[174] = 'h7785;
        exp_re_rom[175] = 'h272ec;
        exp_re_rom[176] = 'h74509;
        exp_re_rom[177] = 'h7ef2407;
        exp_re_rom[178] = 'h7fc2782;
        exp_re_rom[179] = 'h7fe15fb;
        exp_re_rom[180] = 'h7ff4a07;
        exp_re_rom[181] = 'h7fd09ef;
        exp_re_rom[182] = 'h7feb22a;
        exp_re_rom[183] = 'h7feddd9;
        exp_re_rom[184] = 'h7fe03a9;
        exp_re_rom[185] = 'h60fa7;
        exp_re_rom[186] = 'h242e3;
        exp_re_rom[187] = 'h2a0a0;
        exp_re_rom[188] = 'h5390c;
        exp_re_rom[189] = 'h7f478fa;
        exp_re_rom[190] = 'h7fecd1a;
        exp_re_rom[191] = 'heaf7;
        exp_re_rom[192] = 'h4fa4f;
        exp_re_rom[193] = 'h7eb32dc;
        exp_re_rom[194] = 'h7fae141;
        exp_re_rom[195] = 'h7fc639c;
        exp_re_rom[196] = 'h7fbe2a6;
        exp_re_rom[197] = 'h65258;
        exp_re_rom[198] = 'h851b;
        exp_re_rom[199] = 'h59af;
        exp_re_rom[200] = 'h13f3f;
        exp_re_rom[201] = 'h7f8fed4;
        exp_re_rom[202] = 'h7fe5230;
        exp_re_rom[203] = 'h7fedaca;
        exp_re_rom[204] = 'h7ff0ab8;
        exp_re_rom[205] = 'h7ff8b80;
        exp_re_rom[206] = 'h7ff66c6;
        exp_re_rom[207] = 'h7ff76fa;
        exp_re_rom[208] = 'h7ff8e08;
        exp_re_rom[209] = 'h7ff4547;
        exp_re_rom[210] = 'h7ff8f42;
        exp_re_rom[211] = 'h7ffa4e0;
        exp_re_rom[212] = 'h7ffc2be;
        exp_re_rom[213] = 'h7ff2efe;
        exp_re_rom[214] = 'h7ffb89f;
        exp_re_rom[215] = 'h7ffe445;
        exp_re_rom[216] = 'h475c;
        exp_re_rom[217] = 'h7fc5f7e;
        exp_re_rom[218] = 'h7ff6703;
        exp_re_rom[219] = 'h7ffd786;
        exp_re_rom[220] = 'hbfaf;
        exp_re_rom[221] = 'h7f49255;
        exp_re_rom[222] = 'h7fd9a81;
        exp_re_rom[223] = 'h7fdd3d2;
        exp_re_rom[224] = 'h7fccccb;
        exp_re_rom[225] = 'h100d43;
        exp_re_rom[226] = 'h11102;
        exp_re_rom[227] = 'h2398;
        exp_re_rom[228] = 'h7ff7a92;
        exp_re_rom[229] = 'h62474;
        exp_re_rom[230] = 'h8432;
        exp_re_rom[231] = 'h1826;
        exp_re_rom[232] = 'h7ffa2f0;
        exp_re_rom[233] = 'h65664;
        exp_re_rom[234] = 'h8ee4;
        exp_re_rom[235] = 'h1e23;
        exp_re_rom[236] = 'h7ff5f8b;
        exp_re_rom[237] = 'h120203;
        exp_re_rom[238] = 'h22788;
        exp_re_rom[239] = 'h1e92e;
        exp_re_rom[240] = 'h2c039;
        exp_re_rom[241] = 'h7e11df4;
        exp_re_rom[242] = 'h7fefc57;
        exp_re_rom[243] = 'h7fff84f;
        exp_re_rom[244] = 'hc3a2;
        exp_re_rom[245] = 'h7e990f6;
        exp_re_rom[246] = 'h7ff18dc;
        exp_re_rom[247] = 'h7ffad8c;
        exp_re_rom[248] = 'h1c28;
        exp_re_rom[249] = 'h7eef708;
        exp_re_rom[250] = 'h7ff5fc8;
        exp_re_rom[251] = 'h7ffa9a6;
        exp_re_rom[252] = 'h7ffd490;
        exp_re_rom[253] = 'h7f6f934;
        exp_re_rom[254] = 'h7ffc125;
        exp_re_rom[255] = 'h7ffde26;
        exp_re_rom[256] = 'h2;
        exp_re_rom[257] = 'h2f5bce;
        exp_re_rom[258] = 'h7ffab25;
        exp_re_rom[259] = 'h7ffc4f7;
        exp_re_rom[260] = 'h7ffcae3;
        exp_re_rom[261] = 'h7fe9380;
        exp_re_rom[262] = 'h7ffd731;
        exp_re_rom[263] = 'h7ffc759;
        exp_re_rom[264] = 'h7ff98a9;
        exp_re_rom[265] = 'h7f4be0a;
        exp_re_rom[266] = 'h6277;
        exp_re_rom[267] = 'h256e;
        exp_re_rom[268] = 'h7fff82a;
        exp_re_rom[269] = 'h7fb3c6b;
        exp_re_rom[270] = 'h6c32;
        exp_re_rom[271] = 'h4095;
        exp_re_rom[272] = 'h1cdb;
        exp_re_rom[273] = 'h7fd121e;
        exp_re_rom[274] = 'h811a;
        exp_re_rom[275] = 'h59b8;
        exp_re_rom[276] = 'h3267;
        exp_re_rom[277] = 'h7fce0a0;
        exp_re_rom[278] = 'hcc92;
        exp_re_rom[279] = 'ha1d7;
        exp_re_rom[280] = 'h8762;
        exp_re_rom[281] = 'h7fe6cf0;
        exp_re_rom[282] = 'h11b53;
        exp_re_rom[283] = 'h1171f;
        exp_re_rom[284] = 'h14434;
        exp_re_rom[285] = 'h34060;
        exp_re_rom[286] = 'h13ca5;
        exp_re_rom[287] = 'h1ecb9;
        exp_re_rom[288] = 'h379fd;
        exp_re_rom[289] = 'h1bfc67;
        exp_re_rom[290] = 'h7fc5531;
        exp_re_rom[291] = 'h7fea3fa;
        exp_re_rom[292] = 'h7ff932b;
        exp_re_rom[293] = 'h374de;
        exp_re_rom[294] = 'h7fefe07;
        exp_re_rom[295] = 'h7ff980b;
        exp_re_rom[296] = 'h1224;
        exp_re_rom[297] = 'h3c467;
        exp_re_rom[298] = 'h7fef3f9;
        exp_re_rom[299] = 'h7ff813c;
        exp_re_rom[300] = 'h7ffdfe3;
        exp_re_rom[301] = 'h2f23d;
        exp_re_rom[302] = 'h7fe7708;
        exp_re_rom[303] = 'h7fe9211;
        exp_re_rom[304] = 'h7fda400;
        exp_re_rom[305] = 'h7f04781;
        exp_re_rom[306] = 'h496a5;
        exp_re_rom[307] = 'h2d8f0;
        exp_re_rom[308] = 'h319a3;
        exp_re_rom[309] = 'haf16b;
        exp_re_rom[310] = 'h7febe0b;
        exp_re_rom[311] = 'h4f92;
        exp_re_rom[312] = 'h1356b;
        exp_re_rom[313] = 'h63595;
        exp_re_rom[314] = 'h7fef26a;
        exp_re_rom[315] = 'h2940;
        exp_re_rom[316] = 'he7c6;
        exp_re_rom[317] = 'h40dbf;
        exp_re_rom[318] = 'h7fff770;
        exp_re_rom[319] = 'h14e92;
        exp_re_rom[320] = 'h33d4b;
        exp_re_rom[321] = 'h128dfe;
        exp_re_rom[322] = 'h7f9034a;
        exp_re_rom[323] = 'h7fcc923;
        exp_re_rom[324] = 'h7fdc70a;
        exp_re_rom[325] = 'h7fdaf3c;
        exp_re_rom[326] = 'h7ff0ee5;
        exp_re_rom[327] = 'h7ff1d01;
        exp_re_rom[328] = 'h7ff4134;
        exp_re_rom[329] = 'h7ff9bc9;
        exp_re_rom[330] = 'h7ff3da1;
        exp_re_rom[331] = 'h7ff66d7;
        exp_re_rom[332] = 'h7ff854f;
        exp_re_rom[333] = 'h7ffe214;
        exp_re_rom[334] = 'h7ff5fab;
        exp_re_rom[335] = 'h7ff8469;
        exp_re_rom[336] = 'h7ff9325;
        exp_re_rom[337] = 'h7ff8564;
        exp_re_rom[338] = 'h7ffcb4e;
        exp_re_rom[339] = 'h7ffd198;
        exp_re_rom[340] = 'h7ffe98c;
        exp_re_rom[341] = 'h6cb0;
        exp_re_rom[342] = 'h7ff7ce5;
        exp_re_rom[343] = 'h7ffb682;
        exp_re_rom[344] = 'h7ffcafd;
        exp_re_rom[345] = 'h7ffd2f0;
        exp_re_rom[346] = 'h7fff652;
        exp_re_rom[347] = 'hacf;
        exp_re_rom[348] = 'h3cf6;
        exp_re_rom[349] = 'h179be;
        exp_re_rom[350] = 'h7fec2e9;
        exp_re_rom[351] = 'h7ff41cc;
        exp_re_rom[352] = 'h7ff14d6;
        exp_re_rom[353] = 'h7fccffb;
        exp_re_rom[354] = 'h2596d;
        exp_re_rom[355] = 'h149b4;
        exp_re_rom[356] = 'h16208;
        exp_re_rom[357] = 'h34833;
        exp_re_rom[358] = 'h7fec7a6;
        exp_re_rom[359] = 'h7fff978;
        exp_re_rom[360] = 'h6cd8;
        exp_re_rom[361] = 'h17ea5;
        exp_re_rom[362] = 'h7ff83da;
        exp_re_rom[363] = 'h4197;
        exp_re_rom[364] = 'haeb3;
        exp_re_rom[365] = 'h1df0a;
        exp_re_rom[366] = 'h7ffb447;
        exp_re_rom[367] = 'hc245;
        exp_re_rom[368] = 'h1c069;
        exp_re_rom[369] = 'h638a3;
        exp_re_rom[370] = 'h7fafec8;
        exp_re_rom[371] = 'h7fe3508;
        exp_re_rom[372] = 'h7feaef6;
        exp_re_rom[373] = 'h7fcd83d;
        exp_re_rom[374] = 'h41b11;
        exp_re_rom[375] = 'h30631;
        exp_re_rom[376] = 'h465c9;
        exp_re_rom[377] = 'hc99e1;
        exp_re_rom[378] = 'h7f6414c;
        exp_re_rom[379] = 'h7fe07eb;
        exp_re_rom[380] = 'h15639;
        exp_re_rom[381] = 'hbefdb;
        exp_re_rom[382] = 'h7ee1547;
        exp_re_rom[383] = 'h7f74bca;
        exp_re_rom[384] = 'h7f7bfdb;
        exp_re_rom[385] = 'h7f03467;
        exp_re_rom[386] = 'hb1ece;
        exp_re_rom[387] = 'h2dfc0;
        exp_re_rom[388] = 'h1f987;
        exp_re_rom[389] = 'h449eb;
        exp_re_rom[390] = 'h7fae6b3;
        exp_re_rom[391] = 'h7fdf630;
        exp_re_rom[392] = 'h7fe731f;
        exp_re_rom[393] = 'h7fe5e44;
        exp_re_rom[394] = 'h7ff8cf4;
        exp_re_rom[395] = 'h7ff45cd;
        exp_re_rom[396] = 'h7ff4e7e;
        exp_re_rom[397] = 'h7ff7e53;
        exp_re_rom[398] = 'h7ff04bf;
        exp_re_rom[399] = 'h7ff4993;
        exp_re_rom[400] = 'h7ff700f;
        exp_re_rom[401] = 'h7ffd939;
        exp_re_rom[402] = 'h7fe8eb8;
        exp_re_rom[403] = 'h7ff14f9;
        exp_re_rom[404] = 'h7ff0c1a;
        exp_re_rom[405] = 'h7fdf9f9;
        exp_re_rom[406] = 'h3a4c1;
        exp_re_rom[407] = 'h23f99;
        exp_re_rom[408] = 'h39ba4;
        exp_re_rom[409] = 'hb0989;
        exp_re_rom[410] = 'h7ec7caa;
        exp_re_rom[411] = 'h7f97fed;
        exp_re_rom[412] = 'h7fbd274;
        exp_re_rom[413] = 'h7fe1acd;
        exp_re_rom[414] = 'h7f6ce5f;
        exp_re_rom[415] = 'h7f97ee5;
        exp_re_rom[416] = 'h7f863d5;
        exp_re_rom[417] = 'h7f150e7;
        exp_re_rom[418] = 'h11eafb;
        exp_re_rom[419] = 'h2e340;
        exp_re_rom[420] = 'h4e91;
        exp_re_rom[421] = 'h7fe3c82;
        exp_re_rom[422] = 'h28459;
        exp_re_rom[423] = 'h7ff7926;
        exp_re_rom[424] = 'h7fe0d67;
        exp_re_rom[425] = 'h7fa41e2;
        exp_re_rom[426] = 'hb3eb9;
        exp_re_rom[427] = 'h277ed;
        exp_re_rom[428] = 'hd98d;
        exp_re_rom[429] = 'h7ff0530;
        exp_re_rom[430] = 'h59b5f;
        exp_re_rom[431] = 'h1fc9b;
        exp_re_rom[432] = 'h192e5;
        exp_re_rom[433] = 'h2253a;
        exp_re_rom[434] = 'h7fcf944;
        exp_re_rom[435] = 'h7ff657b;
        exp_re_rom[436] = 'h7ff7297;
        exp_re_rom[437] = 'h7fe966c;
        exp_re_rom[438] = 'h4e01c;
        exp_re_rom[439] = 'h1e201;
        exp_re_rom[440] = 'h24e64;
        exp_re_rom[441] = 'h5a641;
        exp_re_rom[442] = 'h7ee0e94;
        exp_re_rom[443] = 'h7fac986;
        exp_re_rom[444] = 'h7fb7687;
        exp_re_rom[445] = 'h7f90305;
        exp_re_rom[446] = 'hcbfe4;
        exp_re_rom[447] = 'h10dc3;
        exp_re_rom[448] = 'h7ff2582;
        exp_re_rom[449] = 'h7fc1e5a;
        exp_re_rom[450] = 'heeb45;
        exp_re_rom[451] = 'h35078;
        exp_re_rom[452] = 'h2206c;
        exp_re_rom[453] = 'h21c1b;
        exp_re_rom[454] = 'h7fdb900;
        exp_re_rom[455] = 'h12bf;
        exp_re_rom[456] = 'h209a;
        exp_re_rom[457] = 'h7ffcf38;
        exp_re_rom[458] = 'h2c387;
        exp_re_rom[459] = 'he253;
        exp_re_rom[460] = 'hc958;
        exp_re_rom[461] = 'h10cd6;
        exp_re_rom[462] = 'h7fde325;
        exp_re_rom[463] = 'h7fff9a1;
        exp_re_rom[464] = 'h2d12;
        exp_re_rom[465] = 'h5663;
        exp_re_rom[466] = 'h7ff5d56;
        exp_re_rom[467] = 'h143a;
        exp_re_rom[468] = 'h1fdd;
        exp_re_rom[469] = 'h7fffa7f;
        exp_re_rom[470] = 'h2d0a8;
        exp_re_rom[471] = 'h1091f;
        exp_re_rom[472] = 'h12e4a;
        exp_re_rom[473] = 'h1e764;
        exp_re_rom[474] = 'h7fa6457;
        exp_re_rom[475] = 'h8545;
        exp_re_rom[476] = 'h1ce3e;
        exp_re_rom[477] = 'h4fa69;
        exp_re_rom[478] = 'h7da065c;
        exp_re_rom[479] = 'h7fae02c;
        exp_re_rom[480] = 'h7fcdd41;
        exp_re_rom[481] = 'h7fd63fb;
        exp_re_rom[482] = 'hf35b;
        exp_re_rom[483] = 'h7fe9de8;
        exp_re_rom[484] = 'h7fe953a;
        exp_re_rom[485] = 'h7fe94bc;
        exp_re_rom[486] = 'h7fe5ffb;
        exp_re_rom[487] = 'h7fe650b;
        exp_re_rom[488] = 'h7fe256a;
        exp_re_rom[489] = 'h7fd5720;
        exp_re_rom[490] = 'he486f;
        exp_re_rom[491] = 'h7ffd2aa;
        exp_re_rom[492] = 'h7feefc0;
        exp_re_rom[493] = 'h7fdd70f;
        exp_re_rom[494] = 'h149330;
        exp_re_rom[495] = 'h77d9;
        exp_re_rom[496] = 'h7ff7614;
        exp_re_rom[497] = 'h7fe575d;
        exp_re_rom[498] = 'h1af462;
        exp_re_rom[499] = 'hef0a;
        exp_re_rom[500] = 'h7fff580;
        exp_re_rom[501] = 'h7ff00ed;
        exp_re_rom[502] = 'h1f7ce0;
        exp_re_rom[503] = 'h12260;
        exp_re_rom[504] = 'h61f5;
        exp_re_rom[505] = 'h7ffd68c;
        exp_re_rom[506] = 'h17511a;
        exp_re_rom[507] = 'ha4ca;
        exp_re_rom[508] = 'h430d;
        exp_re_rom[509] = 'h7fffbbc;
        exp_re_rom[510] = 'h1e93e1;
        exp_re_rom[511] = 'h3f02;
        exp_re_rom[512] = 'h7fffff6;
        exp_re_rom[513] = 'h7ffb0b6;
        exp_re_rom[514] = 'h7c6f83d;
        exp_re_rom[515] = 'h72fc;
        exp_re_rom[516] = 'h21ca;
        exp_re_rom[517] = 'h7ffdade;
        exp_re_rom[518] = 'h7f0ce3f;
        exp_re_rom[519] = 'h7766;
        exp_re_rom[520] = 'h3ca3;
        exp_re_rom[521] = 'h1f7d;
        exp_re_rom[522] = 'h7fef228;
        exp_re_rom[523] = 'h1b7d;
        exp_re_rom[524] = 'h966;
        exp_re_rom[525] = 'h7fff809;
        exp_re_rom[526] = 'h7ff0f1f;
        exp_re_rom[527] = 'h7fff9d1;
        exp_re_rom[528] = 'h7ffe0c5;
        exp_re_rom[529] = 'h7ffb952;
        exp_re_rom[530] = 'h7fc8cf3;
        exp_re_rom[531] = 'h1221;
        exp_re_rom[532] = 'h7ffd237;
        exp_re_rom[533] = 'h7ff81ad;
        exp_re_rom[534] = 'h7fa32bf;
        exp_re_rom[535] = 'h3a44;
        exp_re_rom[536] = 'h7ffa964;
        exp_re_rom[537] = 'h7fecbcb;
        exp_re_rom[538] = 'h7ef6740;
        exp_re_rom[539] = 'h1fac9;
        exp_re_rom[540] = 'h96d2;
        exp_re_rom[541] = 'h7feff4f;
        exp_re_rom[542] = 'h7e40005;
        exp_re_rom[543] = 'h6ee9e;
        exp_re_rom[544] = 'h5d252;
        exp_re_rom[545] = 'h81dd6;
        exp_re_rom[546] = 'h36e16f;
        exp_re_rom[547] = 'h7f94f43;
        exp_re_rom[548] = 'h7fdd170;
        exp_re_rom[549] = 'h7ffb50e;
        exp_re_rom[550] = 'h9232b;
        exp_re_rom[551] = 'h7fdc071;
        exp_re_rom[552] = 'h7ff34c3;
        exp_re_rom[553] = 'h7544;
        exp_re_rom[554] = 'hbb330;
        exp_re_rom[555] = 'h7fc808c;
        exp_re_rom[556] = 'h7fe013c;
        exp_re_rom[557] = 'h7fe8f1f;
        exp_re_rom[558] = 'h7ffcc28;
        exp_re_rom[559] = 'h7fe7f76;
        exp_re_rom[560] = 'h7feb7ce;
        exp_re_rom[561] = 'h7fec0f4;
        exp_re_rom[562] = 'h7fdcf22;
        exp_re_rom[563] = 'h7ff725c;
        exp_re_rom[564] = 'h7ff659f;
        exp_re_rom[565] = 'h7ff9d7a;
        exp_re_rom[566] = 'h25d1d;
        exp_re_rom[567] = 'h7fdfdce;
        exp_re_rom[568] = 'h7fe59ff;
        exp_re_rom[569] = 'h7fe1424;
        exp_re_rom[570] = 'h7f9c996;
        exp_re_rom[571] = 'hf36a;
        exp_re_rom[572] = 'h5305;
        exp_re_rom[573] = 'hded3;
        exp_re_rom[574] = 'h926d9;
        exp_re_rom[575] = 'h7fa9431;
        exp_re_rom[576] = 'h7fbd0a6;
        exp_re_rom[577] = 'h7fa955d;
        exp_re_rom[578] = 'h7ebe1e4;
        exp_re_rom[579] = 'h52d82;
        exp_re_rom[580] = 'h151a5;
        exp_re_rom[581] = 'h7ffe12a;
        exp_re_rom[582] = 'h7fb7a7a;
        exp_re_rom[583] = 'h23023;
        exp_re_rom[584] = 'he6f2;
        exp_re_rom[585] = 'h7046;
        exp_re_rom[586] = 'h7ffbd0e;
        exp_re_rom[587] = 'h77fd;
        exp_re_rom[588] = 'h33f3;
        exp_re_rom[589] = 'h96b;
        exp_re_rom[590] = 'h7ff85e4;
        exp_re_rom[591] = 'h4fd9;
        exp_re_rom[592] = 'h2144;
        exp_re_rom[593] = 'h14ce;
        exp_re_rom[594] = 'h29e8;
        exp_re_rom[595] = 'h7ffef90;
        exp_re_rom[596] = 'h1cb;
        exp_re_rom[597] = 'h2456;
        exp_re_rom[598] = 'h1276c;
        exp_re_rom[599] = 'h7ff14fe;
        exp_re_rom[600] = 'h7ff82ba;
        exp_re_rom[601] = 'h7ffa996;
        exp_re_rom[602] = 'hb06;
        exp_re_rom[603] = 'h7ff7967;
        exp_re_rom[604] = 'h7ffcb0d;
        exp_re_rom[605] = 'h5ae0;
        exp_re_rom[606] = 'h45be6;
        exp_re_rom[607] = 'h7fb12eb;
        exp_re_rom[608] = 'h7fca16b;
        exp_re_rom[609] = 'h7fbf4dc;
        exp_re_rom[610] = 'h7f5070c;
        exp_re_rom[611] = 'h53270;
        exp_re_rom[612] = 'h17c0e;
        exp_re_rom[613] = 'hc634;
        exp_re_rom[614] = 'h192cc;
        exp_re_rom[615] = 'h7fe4b9d;
        exp_re_rom[616] = 'h7feb2be;
        exp_re_rom[617] = 'h7fe650d;
        exp_re_rom[618] = 'h7fcd51d;
        exp_re_rom[619] = 'h7ffb482;
        exp_re_rom[620] = 'h7fe2199;
        exp_re_rom[621] = 'h7fc29ca;
        exp_re_rom[622] = 'h7f1c451;
        exp_re_rom[623] = 'hc266b;
        exp_re_rom[624] = 'h53f33;
        exp_re_rom[625] = 'h46e83;
        exp_re_rom[626] = 'h7e2aa;
        exp_re_rom[627] = 'h7fd1595;
        exp_re_rom[628] = 'h5b83;
        exp_re_rom[629] = 'h2276f;
        exp_re_rom[630] = 'ha36b0;
        exp_re_rom[631] = 'h7f36e52;
        exp_re_rom[632] = 'h7f965a5;
        exp_re_rom[633] = 'h7f9187a;
        exp_re_rom[634] = 'h7f1643c;
        exp_re_rom[635] = 'h835b0;
        exp_re_rom[636] = 'h82f0;
        exp_re_rom[637] = 'h7fd7790;
        exp_re_rom[638] = 'h7f4340f;
        exp_re_rom[639] = 'hdffbc;
        exp_re_rom[640] = 'h58bb1;
        exp_re_rom[641] = 'h45410;
        exp_re_rom[642] = 'h6e329;
        exp_re_rom[643] = 'h7fb516d;
        exp_re_rom[644] = 'h7fe48e7;
        exp_re_rom[645] = 'h7fdbfb7;
        exp_re_rom[646] = 'h7f8b69b;
        exp_re_rom[647] = 'h9b393;
        exp_re_rom[648] = 'h3dadb;
        exp_re_rom[649] = 'h30850;
        exp_re_rom[650] = 'h411fb;
        exp_re_rom[651] = 'h7feae10;
        exp_re_rom[652] = 'h6af6;
        exp_re_rom[653] = 'hadf1;
        exp_re_rom[654] = 'hd9e1;
        exp_re_rom[655] = 'h89f4;
        exp_re_rom[656] = 'hb5ce;
        exp_re_rom[657] = 'hcd9b;
        exp_re_rom[658] = 'h1131c;
        exp_re_rom[659] = 'h4350;
        exp_re_rom[660] = 'hb12b;
        exp_re_rom[661] = 'he9c1;
        exp_re_rom[662] = 'h179e0;
        exp_re_rom[663] = 'h7ffeca7;
        exp_re_rom[664] = 'heb7d;
        exp_re_rom[665] = 'h1a42d;
        exp_re_rom[666] = 'h41944;
        exp_re_rom[667] = 'h7fb09a4;
        exp_re_rom[668] = 'h7ff794a;
        exp_re_rom[669] = 'h124c0;
        exp_re_rom[670] = 'h5ff7a;
        exp_re_rom[671] = 'h7f1b715;
        exp_re_rom[672] = 'h7fa78e5;
        exp_re_rom[673] = 'h7fb219c;
        exp_re_rom[674] = 'h7f84ce2;
        exp_re_rom[675] = 'h840ee;
        exp_re_rom[676] = 'h167ed;
        exp_re_rom[677] = 'h104c7;
        exp_re_rom[678] = 'h3dabb;
        exp_re_rom[679] = 'h7f1dd43;
        exp_re_rom[680] = 'h7f8dbba;
        exp_re_rom[681] = 'h7f77358;
        exp_re_rom[682] = 'h7edbf6b;
        exp_re_rom[683] = 'h2013e9;
        exp_re_rom[684] = 'h6bea3;
        exp_re_rom[685] = 'h26d38;
        exp_re_rom[686] = 'h7fd8a2f;
        exp_re_rom[687] = 'h107e6a;
        exp_re_rom[688] = 'h65ff3;
        exp_re_rom[689] = 'h58b53;
        exp_re_rom[690] = 'h806be;
        exp_re_rom[691] = 'h7f57cb9;
        exp_re_rom[692] = 'h7fef981;
        exp_re_rom[693] = 'h3be7;
        exp_re_rom[694] = 'h187c2;
        exp_re_rom[695] = 'h7fb0f6d;
        exp_re_rom[696] = 'h7fe607d;
        exp_re_rom[697] = 'h7fe2a89;
        exp_re_rom[698] = 'h7fbc293;
        exp_re_rom[699] = 'hc7d30;
        exp_re_rom[700] = 'h2fec6;
        exp_re_rom[701] = 'h1d720;
        exp_re_rom[702] = 'h10fe2;
        exp_re_rom[703] = 'h437bf;
        exp_re_rom[704] = 'h27a71;
        exp_re_rom[705] = 'h2d196;
        exp_re_rom[706] = 'h50beb;
        exp_re_rom[707] = 'h7f34d7e;
        exp_re_rom[708] = 'h7fe036c;
        exp_re_rom[709] = 'h7ff06be;
        exp_re_rom[710] = 'h7ff1551;
        exp_re_rom[711] = 'h229ff;
        exp_re_rom[712] = 'h83b3;
        exp_re_rom[713] = 'h822e;
        exp_re_rom[714] = 'hdb5e;
        exp_re_rom[715] = 'h7fdaad0;
        exp_re_rom[716] = 'h7ffc30c;
        exp_re_rom[717] = 'h7fff85e;
        exp_re_rom[718] = 'h160c;
        exp_re_rom[719] = 'h7ffb3c0;
        exp_re_rom[720] = 'h4c;
        exp_re_rom[721] = 'h6c5;
        exp_re_rom[722] = 'hbe;
        exp_re_rom[723] = 'h65a8;
        exp_re_rom[724] = 'h1d80;
        exp_re_rom[725] = 'h10b4;
        exp_re_rom[726] = 'h7fff317;
        exp_re_rom[727] = 'h12db7;
        exp_re_rom[728] = 'h451c;
        exp_re_rom[729] = 'h2b6e;
        exp_re_rom[730] = 'h58f;
        exp_re_rom[731] = 'h1a5d8;
        exp_re_rom[732] = 'h6b2f;
        exp_re_rom[733] = 'h5055;
        exp_re_rom[734] = 'h2b35;
        exp_re_rom[735] = 'h26294;
        exp_re_rom[736] = 'hca21;
        exp_re_rom[737] = 'hdb9f;
        exp_re_rom[738] = 'h15684;
        exp_re_rom[739] = 'h7f99ab6;
        exp_re_rom[740] = 'h7fff302;
        exp_re_rom[741] = 'h9d18;
        exp_re_rom[742] = 'h1e116;
        exp_re_rom[743] = 'h7eae6de;
        exp_re_rom[744] = 'h7fdc990;
        exp_re_rom[745] = 'h7feaacc;
        exp_re_rom[746] = 'h7ff1880;
        exp_re_rom[747] = 'h7f968f1;
        exp_re_rom[748] = 'h7fdef95;
        exp_re_rom[749] = 'h7fd7409;
        exp_re_rom[750] = 'h7fb389c;
        exp_re_rom[751] = 'h3fb7b8;
        exp_re_rom[752] = 'h3ebe7;
        exp_re_rom[753] = 'h20baa;
        exp_re_rom[754] = 'h16be7;
        exp_re_rom[755] = 'h17b9d;
        exp_re_rom[756] = 'h10c8a;
        exp_re_rom[757] = 'h10892;
        exp_re_rom[758] = 'h144ca;
        exp_re_rom[759] = 'h7f06a50;
        exp_re_rom[760] = 'h16fe;
        exp_re_rom[761] = 'h6b94;
        exp_re_rom[762] = 'hc392;
        exp_re_rom[763] = 'h7e5513a;
        exp_re_rom[764] = 'h7ffc508;
        exp_re_rom[765] = 'h107e;
        exp_re_rom[766] = 'h3fc9;
        exp_re_rom[767] = 'h7d31140;
        exp_re_rom[768] = 'h7fffff2;
        exp_re_rom[769] = 'h265e;
        exp_re_rom[770] = 'h535f;
        exp_re_rom[771] = 'h16bf0f;
        exp_re_rom[772] = 'h7ffda8d;
        exp_re_rom[773] = 'h8d6;
        exp_re_rom[774] = 'h323b;
        exp_re_rom[775] = 'h8a2b5;
        exp_re_rom[776] = 'h7ffc109;
        exp_re_rom[777] = 'h7ffe080;
        exp_re_rom[778] = 'h7ffe471;
        exp_re_rom[779] = 'h7fe6806;
        exp_re_rom[780] = 'h103e;
        exp_re_rom[781] = 'h701;
        exp_re_rom[782] = 'h7fffcc8;
        exp_re_rom[783] = 'h7fe8f41;
        exp_re_rom[784] = 'h2e4b;
        exp_re_rom[785] = 'h24e8;
        exp_re_rom[786] = 'h263c;
        exp_re_rom[787] = 'h6cb0;
        exp_re_rom[788] = 'h21c5;
        exp_re_rom[789] = 'h2e1c;
        exp_re_rom[790] = 'h475c;
        exp_re_rom[791] = 'h23f47;
        exp_re_rom[792] = 'h7fff050;
        exp_re_rom[793] = 'h1956;
        exp_re_rom[794] = 'h41e9;
        exp_re_rom[795] = 'h25f15;
        exp_re_rom[796] = 'h7ffe3e8;
        exp_re_rom[797] = 'h2c36;
        exp_re_rom[798] = 'ha239;
        exp_re_rom[799] = 'h8892b;
        exp_re_rom[800] = 'h7fe4d8f;
        exp_re_rom[801] = 'h7fec13b;
        exp_re_rom[802] = 'h7fe5a87;
        exp_re_rom[803] = 'h7f4c75c;
        exp_re_rom[804] = 'h1a493;
        exp_re_rom[805] = 'hc3e2;
        exp_re_rom[806] = 'h8235;
        exp_re_rom[807] = 'h7ff6fa5;
        exp_re_rom[808] = 'h10426;
        exp_re_rom[809] = 'h13699;
        exp_re_rom[810] = 'h2165b;
        exp_re_rom[811] = 'hd5e86;
        exp_re_rom[812] = 'h7fddbb1;
        exp_re_rom[813] = 'h7ffde9d;
        exp_re_rom[814] = 'h2226a;
        exp_re_rom[815] = 'h1b718b;
        exp_re_rom[816] = 'h7f5bc12;
        exp_re_rom[817] = 'h7f83e5b;
        exp_re_rom[818] = 'h7f5e89f;
        exp_re_rom[819] = 'h7d0ebdc;
        exp_re_rom[820] = 'h93f53;
        exp_re_rom[821] = 'h2edbd;
        exp_re_rom[822] = 'h8c99;
        exp_re_rom[823] = 'h7f87112;
        exp_re_rom[824] = 'h34a17;
        exp_re_rom[825] = 'h17dbd;
        exp_re_rom[826] = 'h811e;
        exp_re_rom[827] = 'h7fc7302;
        exp_re_rom[828] = 'h1f610;
        exp_re_rom[829] = 'hb3fd;
        exp_re_rom[830] = 'h7ff5acc;
        exp_re_rom[831] = 'h7f4d760;
        exp_re_rom[832] = 'h66901;
        exp_re_rom[833] = 'h462e2;
        exp_re_rom[834] = 'h4f698;
        exp_re_rom[835] = 'hfc545;
        exp_re_rom[836] = 'h7fc8054;
        exp_re_rom[837] = 'h7ff503a;
        exp_re_rom[838] = 'h2c01;
        exp_re_rom[839] = 'h1f879;
        exp_re_rom[840] = 'h7ff735a;
        exp_re_rom[841] = 'h7fffecd;
        exp_re_rom[842] = 'h3bbd;
        exp_re_rom[843] = 'hdbbd;
        exp_re_rom[844] = 'h7fff1d5;
        exp_re_rom[845] = 'h29c8;
        exp_re_rom[846] = 'h43df;
        exp_re_rom[847] = 'h8795;
        exp_re_rom[848] = 'h1f5d;
        exp_re_rom[849] = 'h3222;
        exp_re_rom[850] = 'h2242;
        exp_re_rom[851] = 'h7ff387a;
        exp_re_rom[852] = 'h1488a;
        exp_re_rom[853] = 'h1151a;
        exp_re_rom[854] = 'h165dd;
        exp_re_rom[855] = 'h40c7a;
        exp_re_rom[856] = 'h7fe9941;
        exp_re_rom[857] = 'h7ffb406;
        exp_re_rom[858] = 'h7ffe4fc;
        exp_re_rom[859] = 'h7ff06ed;
        exp_re_rom[860] = 'h1ad2e;
        exp_re_rom[861] = 'h199b2;
        exp_re_rom[862] = 'h27717;
        exp_re_rom[863] = 'h87414;
        exp_re_rom[864] = 'h7fb6858;
        exp_re_rom[865] = 'h7fe8b09;
        exp_re_rom[866] = 'h7ffaa83;
        exp_re_rom[867] = 'h2dd12;
        exp_re_rom[868] = 'h7fc199c;
        exp_re_rom[869] = 'h7fd8a1d;
        exp_re_rom[870] = 'h7fd426c;
        exp_re_rom[871] = 'h7f91b46;
        exp_re_rom[872] = 'h380fe;
        exp_re_rom[873] = 'hefaf;
        exp_re_rom[874] = 'h3e00;
        exp_re_rom[875] = 'h7fef8f9;
        exp_re_rom[876] = 'h18c4d;
        exp_re_rom[877] = 'hd288;
        exp_re_rom[878] = 'haa93;
        exp_re_rom[879] = 'h71a3;
        exp_re_rom[880] = 'h15129;
        exp_re_rom[881] = 'h19c75;
        exp_re_rom[882] = 'h2f9d0;
        exp_re_rom[883] = 'hbe3d2;
        exp_re_rom[884] = 'h7f24088;
        exp_re_rom[885] = 'h7f80873;
        exp_re_rom[886] = 'h7f602e9;
        exp_re_rom[887] = 'h7e3136f;
        exp_re_rom[888] = 'h1a61ed;
        exp_re_rom[889] = 'ha8357;
        exp_re_rom[890] = 'h8190e;
        exp_re_rom[891] = 'h9fb93;
        exp_re_rom[892] = 'h264ef;
        exp_re_rom[893] = 'h612a3;
        exp_re_rom[894] = 'ha4469;
        exp_re_rom[895] = 'h1eb562;
        exp_re_rom[896] = 'h7e0f4cf;
        exp_re_rom[897] = 'h7f4dc59;
        exp_re_rom[898] = 'h7f7e5ca;
        exp_re_rom[899] = 'h7f49b20;
        exp_re_rom[900] = 'h5512d;
        exp_re_rom[901] = 'h9c0f;
        exp_re_rom[902] = 'h435b;
        exp_re_rom[903] = 'h19bde;
        exp_re_rom[904] = 'h7fcb4cf;
        exp_re_rom[905] = 'h7fe840a;
        exp_re_rom[906] = 'h7fefcca;
        exp_re_rom[907] = 'h7ffbb63;
        exp_re_rom[908] = 'h7fdd4f0;
        exp_re_rom[909] = 'h7fea631;
        exp_re_rom[910] = 'h7fedbab;
        exp_re_rom[911] = 'h7ff188d;
        exp_re_rom[912] = 'h7fe95bd;
        exp_re_rom[913] = 'h7fed637;
        exp_re_rom[914] = 'h7feed74;
        exp_re_rom[915] = 'h7ff3a3b;
        exp_re_rom[916] = 'h7fde8e6;
        exp_re_rom[917] = 'h7fe433b;
        exp_re_rom[918] = 'h7fe07ed;
        exp_re_rom[919] = 'h7fcd167;
        exp_re_rom[920] = 'h1439c;
        exp_re_rom[921] = 'h7ff24d7;
        exp_re_rom[922] = 'h7fe6250;
        exp_re_rom[923] = 'h7fc94af;
        exp_re_rom[924] = 'h2b164;
        exp_re_rom[925] = 'h7ff872b;
        exp_re_rom[926] = 'h7fe493b;
        exp_re_rom[927] = 'h7fae891;
        exp_re_rom[928] = 'h87081;
        exp_re_rom[929] = 'h2331d;
        exp_re_rom[930] = 'h1442d;
        exp_re_rom[931] = 'h17f42;
        exp_re_rom[932] = 'h7fd51a9;
        exp_re_rom[933] = 'h7fe7dba;
        exp_re_rom[934] = 'h7fdbbdd;
        exp_re_rom[935] = 'h7fa0564;
        exp_re_rom[936] = 'hc1cb5;
        exp_re_rom[937] = 'h368c4;
        exp_re_rom[938] = 'h25db7;
        exp_re_rom[939] = 'h31bf3;
        exp_re_rom[940] = 'h7fb6d89;
        exp_re_rom[941] = 'h7fe75ce;
        exp_re_rom[942] = 'h7fdef9d;
        exp_re_rom[943] = 'h7fa5bcb;
        exp_re_rom[944] = 'hebc87;
        exp_re_rom[945] = 'h46408;
        exp_re_rom[946] = 'h36d18;
        exp_re_rom[947] = 'h4c1e5;
        exp_re_rom[948] = 'h7f8eff9;
        exp_re_rom[949] = 'h7fe8daa;
        exp_re_rom[950] = 'h7fe5f14;
        exp_re_rom[951] = 'h7fada91;
        exp_re_rom[952] = 'h1429ae;
        exp_re_rom[953] = 'h745b7;
        exp_re_rom[954] = 'h783ba;
        exp_re_rom[955] = 'he0f56;
        exp_re_rom[956] = 'h7def96f;
        exp_re_rom[957] = 'h7f9e569;
        exp_re_rom[958] = 'h7fd21d0;
        exp_re_rom[959] = 'h7ff2fc7;
        exp_re_rom[960] = 'h7f84e7e;
        exp_re_rom[961] = 'h7fcb7c8;
        exp_re_rom[962] = 'h7fcd383;
        exp_re_rom[963] = 'h7fb09c2;
        exp_re_rom[964] = 'hb0d76;
        exp_re_rom[965] = 'h15d2b;
        exp_re_rom[966] = 'h5f94;
        exp_re_rom[967] = 'h7ffdccb;
        exp_re_rom[968] = 'h11e34;
        exp_re_rom[969] = 'h11aa;
        exp_re_rom[970] = 'h7ffd09f;
        exp_re_rom[971] = 'h7ff563b;
        exp_re_rom[972] = 'h2fbbc;
        exp_re_rom[973] = 'h87cc;
        exp_re_rom[974] = 'h4bc1;
        exp_re_rom[975] = 'h36a9;
        exp_re_rom[976] = 'h1fd6;
        exp_re_rom[977] = 'h2601;
        exp_re_rom[978] = 'h2de2;
        exp_re_rom[979] = 'h55fa;
        exp_re_rom[980] = 'h7fe89f9;
        exp_re_rom[981] = 'h7ffcf0f;
        exp_re_rom[982] = 'h7ffefca;
        exp_re_rom[983] = 'h1639;
        exp_re_rom[984] = 'h7fecb82;
        exp_re_rom[985] = 'h7ffcf0c;
        exp_re_rom[986] = 'h7ffff6f;
        exp_re_rom[987] = 'h7f85;
        exp_re_rom[988] = 'h7f9619c;
        exp_re_rom[989] = 'h7fe8999;
        exp_re_rom[990] = 'h7fe976a;
        exp_re_rom[991] = 'h7fdc1ba;
        exp_re_rom[992] = 'hbfe9f;
        exp_re_rom[993] = 'hfbd7;
        exp_re_rom[994] = 'h50eb;
        exp_re_rom[995] = 'h7fffd5e;
        exp_re_rom[996] = 'h161aa;
        exp_re_rom[997] = 'haa0;
        exp_re_rom[998] = 'h7ffd72d;
        exp_re_rom[999] = 'h7ff8009;
        exp_re_rom[1000] = 'h50f42;
        exp_re_rom[1001] = 'h6008;
        exp_re_rom[1002] = 'h1f69;
        exp_re_rom[1003] = 'h7fffe1e;
        exp_re_rom[1004] = 'h3530;
        exp_re_rom[1005] = 'h7ffd7d9;
        exp_re_rom[1006] = 'h7ffac3c;
        exp_re_rom[1007] = 'h7ff3cbd;
        exp_re_rom[1008] = 'hbaf20;
        exp_re_rom[1009] = 'ha5e9;
        exp_re_rom[1010] = 'h447c;
        exp_re_rom[1011] = 'hc3e;
        exp_re_rom[1012] = 'h386ec;
        exp_re_rom[1013] = 'h39c3;
        exp_re_rom[1014] = 'h15be;
        exp_re_rom[1015] = 'h7ffef6c;
        exp_re_rom[1016] = 'h5ff0d;
        exp_re_rom[1017] = 'h3d58;
        exp_re_rom[1018] = 'h1f68;
        exp_re_rom[1019] = 'hd52;
        exp_re_rom[1020] = 'h2d027;
        exp_re_rom[1021] = 'h155a;
        exp_re_rom[1022] = 'haed;
        exp_re_rom[1023] = 'h4c0;
    end
    else begin
        exp_re_rom[0] = 'h7fffeda;
        exp_re_rom[1] = 'h4d3;
        exp_re_rom[2] = 'hb00;
        exp_re_rom[3] = 'h1569;
        exp_re_rom[4] = 'h2d02f;
        exp_re_rom[5] = 'hd71;
        exp_re_rom[6] = 'h1f74;
        exp_re_rom[7] = 'h3d69;
        exp_re_rom[8] = 'h5ff03;
        exp_re_rom[9] = 'h7ffef5f;
        exp_re_rom[10] = 'h15cb;
        exp_re_rom[11] = 'h39b9;
        exp_re_rom[12] = 'h386ed;
        exp_re_rom[13] = 'hc31;
        exp_re_rom[14] = 'h449a;
        exp_re_rom[15] = 'ha615;
        exp_re_rom[16] = 'hbaf1b;
        exp_re_rom[17] = 'h7ff3ce6;
        exp_re_rom[18] = 'h7ffac3f;
        exp_re_rom[19] = 'h7ffd7c1;
        exp_re_rom[20] = 'h352e;
        exp_re_rom[21] = 'h7fffe2e;
        exp_re_rom[22] = 'h1f6c;
        exp_re_rom[23] = 'h6008;
        exp_re_rom[24] = 'h50f46;
        exp_re_rom[25] = 'h7ff8019;
        exp_re_rom[26] = 'h7ffd729;
        exp_re_rom[27] = 'ha99;
        exp_re_rom[28] = 'h161a8;
        exp_re_rom[29] = 'h7fffd5c;
        exp_re_rom[30] = 'h50de;
        exp_re_rom[31] = 'hfbd3;
        exp_re_rom[32] = 'hbfe99;
        exp_re_rom[33] = 'h7fdc1b0;
        exp_re_rom[34] = 'h7fe9761;
        exp_re_rom[35] = 'h7fe89b2;
        exp_re_rom[36] = 'h7f9619d;
        exp_re_rom[37] = 'h7f74;
        exp_re_rom[38] = 'h7ffff65;
        exp_re_rom[39] = 'h7ffcf03;
        exp_re_rom[40] = 'h7fecb90;
        exp_re_rom[41] = 'h1626;
        exp_re_rom[42] = 'h7ffefca;
        exp_re_rom[43] = 'h7ffcf05;
        exp_re_rom[44] = 'h7fe89ef;
        exp_re_rom[45] = 'h55f2;
        exp_re_rom[46] = 'h2ddd;
        exp_re_rom[47] = 'h260a;
        exp_re_rom[48] = 'h1fd6;
        exp_re_rom[49] = 'h36a2;
        exp_re_rom[50] = 'h4bc8;
        exp_re_rom[51] = 'h87d2;
        exp_re_rom[52] = 'h2fbb7;
        exp_re_rom[53] = 'h7ff5622;
        exp_re_rom[54] = 'h7ffd0af;
        exp_re_rom[55] = 'h11a5;
        exp_re_rom[56] = 'h11e38;
        exp_re_rom[57] = 'h7ffdcb8;
        exp_re_rom[58] = 'h5f9a;
        exp_re_rom[59] = 'h15d22;
        exp_re_rom[60] = 'hb0d81;
        exp_re_rom[61] = 'h7fb09ce;
        exp_re_rom[62] = 'h7fcd384;
        exp_re_rom[63] = 'h7fcb7c9;
        exp_re_rom[64] = 'h7f84e7e;
        exp_re_rom[65] = 'h7ff2fc4;
        exp_re_rom[66] = 'h7fd21bf;
        exp_re_rom[67] = 'h7f9e571;
        exp_re_rom[68] = 'h7def95c;
        exp_re_rom[69] = 'he0f6a;
        exp_re_rom[70] = 'h783c7;
        exp_re_rom[71] = 'h745c3;
        exp_re_rom[72] = 'h1429aa;
        exp_re_rom[73] = 'h7fada95;
        exp_re_rom[74] = 'h7fe5ef8;
        exp_re_rom[75] = 'h7fe8dc1;
        exp_re_rom[76] = 'h7f8eff8;
        exp_re_rom[77] = 'h4c1c6;
        exp_re_rom[78] = 'h36d11;
        exp_re_rom[79] = 'h46405;
        exp_re_rom[80] = 'hebc95;
        exp_re_rom[81] = 'h7fa5c08;
        exp_re_rom[82] = 'h7fdef7b;
        exp_re_rom[83] = 'h7fe75c6;
        exp_re_rom[84] = 'h7fb6d8c;
        exp_re_rom[85] = 'h31c2a;
        exp_re_rom[86] = 'h25d91;
        exp_re_rom[87] = 'h368c1;
        exp_re_rom[88] = 'hc1cb5;
        exp_re_rom[89] = 'h7fa0559;
        exp_re_rom[90] = 'h7fdbbd2;
        exp_re_rom[91] = 'h7fe7db9;
        exp_re_rom[92] = 'h7fd51b4;
        exp_re_rom[93] = 'h17f47;
        exp_re_rom[94] = 'h143e9;
        exp_re_rom[95] = 'h23312;
        exp_re_rom[96] = 'h8708d;
        exp_re_rom[97] = 'h7fae883;
        exp_re_rom[98] = 'h7fe4944;
        exp_re_rom[99] = 'h7ff872a;
        exp_re_rom[100] = 'h2b16c;
        exp_re_rom[101] = 'h7fc94c6;
        exp_re_rom[102] = 'h7fe6270;
        exp_re_rom[103] = 'h7ff24b7;
        exp_re_rom[104] = 'h1439e;
        exp_re_rom[105] = 'h7fcd156;
        exp_re_rom[106] = 'h7fe07df;
        exp_re_rom[107] = 'h7fe433a;
        exp_re_rom[108] = 'h7fde8e0;
        exp_re_rom[109] = 'h7ff3a2e;
        exp_re_rom[110] = 'h7feed68;
        exp_re_rom[111] = 'h7fed630;
        exp_re_rom[112] = 'h7fe95bc;
        exp_re_rom[113] = 'h7ff18a2;
        exp_re_rom[114] = 'h7fedbb5;
        exp_re_rom[115] = 'h7fea64c;
        exp_re_rom[116] = 'h7fdd4ef;
        exp_re_rom[117] = 'h7ffbb4f;
        exp_re_rom[118] = 'h7fefcc9;
        exp_re_rom[119] = 'h7fe840e;
        exp_re_rom[120] = 'h7fcb4dc;
        exp_re_rom[121] = 'h19bd8;
        exp_re_rom[122] = 'h4353;
        exp_re_rom[123] = 'h9c1a;
        exp_re_rom[124] = 'h55128;
        exp_re_rom[125] = 'h7f49b1a;
        exp_re_rom[126] = 'h7f7e5b5;
        exp_re_rom[127] = 'h7f4dc4d;
        exp_re_rom[128] = 'h7e0f4cf;
        exp_re_rom[129] = 'h1eb536;
        exp_re_rom[130] = 'ha444d;
        exp_re_rom[131] = 'h612ac;
        exp_re_rom[132] = 'h264f9;
        exp_re_rom[133] = 'h9fb95;
        exp_re_rom[134] = 'h81904;
        exp_re_rom[135] = 'ha8352;
        exp_re_rom[136] = 'h1a61e1;
        exp_re_rom[137] = 'h7e3137e;
        exp_re_rom[138] = 'h7f6030a;
        exp_re_rom[139] = 'h7f80874;
        exp_re_rom[140] = 'h7f2408b;
        exp_re_rom[141] = 'hbe3d0;
        exp_re_rom[142] = 'h2f9e8;
        exp_re_rom[143] = 'h19c75;
        exp_re_rom[144] = 'h15122;
        exp_re_rom[145] = 'h71bc;
        exp_re_rom[146] = 'haa6e;
        exp_re_rom[147] = 'hd283;
        exp_re_rom[148] = 'h18c4b;
        exp_re_rom[149] = 'h7fef902;
        exp_re_rom[150] = 'h3de6;
        exp_re_rom[151] = 'hefbc;
        exp_re_rom[152] = 'h380fe;
        exp_re_rom[153] = 'h7f91b54;
        exp_re_rom[154] = 'h7fd4280;
        exp_re_rom[155] = 'h7fd8a30;
        exp_re_rom[156] = 'h7fc19a6;
        exp_re_rom[157] = 'h2dd19;
        exp_re_rom[158] = 'h7ffaaa2;
        exp_re_rom[159] = 'h7fe8b03;
        exp_re_rom[160] = 'h7fb684c;
        exp_re_rom[161] = 'h873fc;
        exp_re_rom[162] = 'h27710;
        exp_re_rom[163] = 'h1999d;
        exp_re_rom[164] = 'h1ad2e;
        exp_re_rom[165] = 'h7ff06ea;
        exp_re_rom[166] = 'h7ffe4ec;
        exp_re_rom[167] = 'h7ffb402;
        exp_re_rom[168] = 'h7fe9942;
        exp_re_rom[169] = 'h40c76;
        exp_re_rom[170] = 'h165db;
        exp_re_rom[171] = 'h1151d;
        exp_re_rom[172] = 'h14882;
        exp_re_rom[173] = 'h7ff387a;
        exp_re_rom[174] = 'h223c;
        exp_re_rom[175] = 'h321b;
        exp_re_rom[176] = 'h1f5d;
        exp_re_rom[177] = 'h879d;
        exp_re_rom[178] = 'h43d9;
        exp_re_rom[179] = 'h29ce;
        exp_re_rom[180] = 'h7fff1d7;
        exp_re_rom[181] = 'hdbc1;
        exp_re_rom[182] = 'h3bcd;
        exp_re_rom[183] = 'h7fffec7;
        exp_re_rom[184] = 'h7ff735c;
        exp_re_rom[185] = 'h1f86c;
        exp_re_rom[186] = 'h2bf8;
        exp_re_rom[187] = 'h7ff503b;
        exp_re_rom[188] = 'h7fc804e;
        exp_re_rom[189] = 'hfc53f;
        exp_re_rom[190] = 'h4f688;
        exp_re_rom[191] = 'h4630c;
        exp_re_rom[192] = 'h66901;
        exp_re_rom[193] = 'h7f4d761;
        exp_re_rom[194] = 'h7ff5ac9;
        exp_re_rom[195] = 'hb3e9;
        exp_re_rom[196] = 'h1f601;
        exp_re_rom[197] = 'h7fc730e;
        exp_re_rom[198] = 'h8116;
        exp_re_rom[199] = 'h17db6;
        exp_re_rom[200] = 'h34a0d;
        exp_re_rom[201] = 'h7f8711a;
        exp_re_rom[202] = 'h8ca1;
        exp_re_rom[203] = 'h2edbe;
        exp_re_rom[204] = 'h93f4f;
        exp_re_rom[205] = 'h7d0ebd8;
        exp_re_rom[206] = 'h7f5e8a4;
        exp_re_rom[207] = 'h7f83e60;
        exp_re_rom[208] = 'h7f5bc0e;
        exp_re_rom[209] = 'h1b718b;
        exp_re_rom[210] = 'h22260;
        exp_re_rom[211] = 'h7ffde9a;
        exp_re_rom[212] = 'h7fddbb3;
        exp_re_rom[213] = 'hd5e8b;
        exp_re_rom[214] = 'h21645;
        exp_re_rom[215] = 'h1369c;
        exp_re_rom[216] = 'h1041e;
        exp_re_rom[217] = 'h7ff6fc0;
        exp_re_rom[218] = 'h8240;
        exp_re_rom[219] = 'hc3ec;
        exp_re_rom[220] = 'h1a49b;
        exp_re_rom[221] = 'h7f4c75b;
        exp_re_rom[222] = 'h7fe5abb;
        exp_re_rom[223] = 'h7fec13a;
        exp_re_rom[224] = 'h7fe4d8f;
        exp_re_rom[225] = 'h88923;
        exp_re_rom[226] = 'ha233;
        exp_re_rom[227] = 'h2c2d;
        exp_re_rom[228] = 'h7ffe3e7;
        exp_re_rom[229] = 'h25efe;
        exp_re_rom[230] = 'h41c7;
        exp_re_rom[231] = 'h1969;
        exp_re_rom[232] = 'h7fff043;
        exp_re_rom[233] = 'h23f4c;
        exp_re_rom[234] = 'h4773;
        exp_re_rom[235] = 'h2e1c;
        exp_re_rom[236] = 'h21c2;
        exp_re_rom[237] = 'h6ca9;
        exp_re_rom[238] = 'h2655;
        exp_re_rom[239] = 'h24d6;
        exp_re_rom[240] = 'h2e4c;
        exp_re_rom[241] = 'h7fe8f3d;
        exp_re_rom[242] = 'h7fffcb5;
        exp_re_rom[243] = 'h715;
        exp_re_rom[244] = 'h1043;
        exp_re_rom[245] = 'h7fe680c;
        exp_re_rom[246] = 'h7ffe476;
        exp_re_rom[247] = 'h7ffe08a;
        exp_re_rom[248] = 'h7ffc107;
        exp_re_rom[249] = 'h8a2a1;
        exp_re_rom[250] = 'h3233;
        exp_re_rom[251] = 'h8d8;
        exp_re_rom[252] = 'h7ffda8f;
        exp_re_rom[253] = 'h16bf25;
        exp_re_rom[254] = 'h535b;
        exp_re_rom[255] = 'h2655;
        exp_re_rom[256] = 'h7fffff2;
        exp_re_rom[257] = 'h7d3114d;
        exp_re_rom[258] = 'h3fb2;
        exp_re_rom[259] = 'h108e;
        exp_re_rom[260] = 'h7ffc506;
        exp_re_rom[261] = 'h7e55136;
        exp_re_rom[262] = 'hc381;
        exp_re_rom[263] = 'h6b88;
        exp_re_rom[264] = 'h1709;
        exp_re_rom[265] = 'h7f06a63;
        exp_re_rom[266] = 'h144ab;
        exp_re_rom[267] = 'h1086a;
        exp_re_rom[268] = 'h10c8b;
        exp_re_rom[269] = 'h17ba8;
        exp_re_rom[270] = 'h16bd3;
        exp_re_rom[271] = 'h20ba2;
        exp_re_rom[272] = 'h3ebeb;
        exp_re_rom[273] = 'h3fb7a1;
        exp_re_rom[274] = 'h7fb38aa;
        exp_re_rom[275] = 'h7fd73fd;
        exp_re_rom[276] = 'h7fdef91;
        exp_re_rom[277] = 'h7f968fd;
        exp_re_rom[278] = 'h7ff1882;
        exp_re_rom[279] = 'h7feaad2;
        exp_re_rom[280] = 'h7fdc992;
        exp_re_rom[281] = 'h7eae6d6;
        exp_re_rom[282] = 'h1e125;
        exp_re_rom[283] = 'h9d25;
        exp_re_rom[284] = 'h7fff300;
        exp_re_rom[285] = 'h7f99abb;
        exp_re_rom[286] = 'h156a3;
        exp_re_rom[287] = 'hdbb5;
        exp_re_rom[288] = 'hca16;
        exp_re_rom[289] = 'h2628f;
        exp_re_rom[290] = 'h2b4f;
        exp_re_rom[291] = 'h505b;
        exp_re_rom[292] = 'h6b3a;
        exp_re_rom[293] = 'h1a5e4;
        exp_re_rom[294] = 'h5a4;
        exp_re_rom[295] = 'h2b61;
        exp_re_rom[296] = 'h4513;
        exp_re_rom[297] = 'h12da8;
        exp_re_rom[298] = 'h7fff319;
        exp_re_rom[299] = 'h10b5;
        exp_re_rom[300] = 'h1d91;
        exp_re_rom[301] = 'h65a6;
        exp_re_rom[302] = 'hc1;
        exp_re_rom[303] = 'h6d7;
        exp_re_rom[304] = 'h4a;
        exp_re_rom[305] = 'h7ffb3be;
        exp_re_rom[306] = 'h1601;
        exp_re_rom[307] = 'h7fff85b;
        exp_re_rom[308] = 'h7ffc313;
        exp_re_rom[309] = 'h7fdaacd;
        exp_re_rom[310] = 'hdb45;
        exp_re_rom[311] = 'h821f;
        exp_re_rom[312] = 'h83b3;
        exp_re_rom[313] = 'h22a00;
        exp_re_rom[314] = 'h7ff1554;
        exp_re_rom[315] = 'h7ff06b6;
        exp_re_rom[316] = 'h7fe035f;
        exp_re_rom[317] = 'h7f34d76;
        exp_re_rom[318] = 'h50be1;
        exp_re_rom[319] = 'h2d189;
        exp_re_rom[320] = 'h27a71;
        exp_re_rom[321] = 'h437c6;
        exp_re_rom[322] = 'h11002;
        exp_re_rom[323] = 'h1d741;
        exp_re_rom[324] = 'h2feb2;
        exp_re_rom[325] = 'hc7d38;
        exp_re_rom[326] = 'h7fbc29d;
        exp_re_rom[327] = 'h7fe2a74;
        exp_re_rom[328] = 'h7fe6094;
        exp_re_rom[329] = 'h7fb0f5b;
        exp_re_rom[330] = 'h187d2;
        exp_re_rom[331] = 'h3bf4;
        exp_re_rom[332] = 'h7fef982;
        exp_re_rom[333] = 'h7f57cb7;
        exp_re_rom[334] = 'h806e0;
        exp_re_rom[335] = 'h58b6d;
        exp_re_rom[336] = 'h65fed;
        exp_re_rom[337] = 'h107e55;
        exp_re_rom[338] = 'h7fd8a43;
        exp_re_rom[339] = 'h26d22;
        exp_re_rom[340] = 'h6bea9;
        exp_re_rom[341] = 'h2013f8;
        exp_re_rom[342] = 'h7edbf67;
        exp_re_rom[343] = 'h7f77356;
        exp_re_rom[344] = 'h7f8dbbf;
        exp_re_rom[345] = 'h7f1dd51;
        exp_re_rom[346] = 'h3dabe;
        exp_re_rom[347] = 'h104c5;
        exp_re_rom[348] = 'h167e4;
        exp_re_rom[349] = 'h840f8;
        exp_re_rom[350] = 'h7f84cf7;
        exp_re_rom[351] = 'h7fb2189;
        exp_re_rom[352] = 'h7fa78ce;
        exp_re_rom[353] = 'h7f1b6e4;
        exp_re_rom[354] = 'h5ff62;
        exp_re_rom[355] = 'h124c8;
        exp_re_rom[356] = 'h7ff7940;
        exp_re_rom[357] = 'h7fb0984;
        exp_re_rom[358] = 'h4193d;
        exp_re_rom[359] = 'h1a42f;
        exp_re_rom[360] = 'heb74;
        exp_re_rom[361] = 'h7ffecaf;
        exp_re_rom[362] = 'h179e8;
        exp_re_rom[363] = 'he9b8;
        exp_re_rom[364] = 'hb128;
        exp_re_rom[365] = 'h435a;
        exp_re_rom[366] = 'h11309;
        exp_re_rom[367] = 'hcd9d;
        exp_re_rom[368] = 'hb5cc;
        exp_re_rom[369] = 'h8a16;
        exp_re_rom[370] = 'hd9f2;
        exp_re_rom[371] = 'haddd;
        exp_re_rom[372] = 'h6aec;
        exp_re_rom[373] = 'h7feae2b;
        exp_re_rom[374] = 'h411df;
        exp_re_rom[375] = 'h3086a;
        exp_re_rom[376] = 'h3dac0;
        exp_re_rom[377] = 'h9b38c;
        exp_re_rom[378] = 'h7f8b6af;
        exp_re_rom[379] = 'h7fdbfb0;
        exp_re_rom[380] = 'h7fe48fb;
        exp_re_rom[381] = 'h7fb5170;
        exp_re_rom[382] = 'h6e351;
        exp_re_rom[383] = 'h4540f;
        exp_re_rom[384] = 'h58bb1;
        exp_re_rom[385] = 'hdffa0;
        exp_re_rom[386] = 'h7f43425;
        exp_re_rom[387] = 'h7fd779d;
        exp_re_rom[388] = 'h82f2;
        exp_re_rom[389] = 'h835a9;
        exp_re_rom[390] = 'h7f1645a;
        exp_re_rom[391] = 'h7f9188e;
        exp_re_rom[392] = 'h7f9658c;
        exp_re_rom[393] = 'h7f36e54;
        exp_re_rom[394] = 'ha369a;
        exp_re_rom[395] = 'h22767;
        exp_re_rom[396] = 'h5b86;
        exp_re_rom[397] = 'h7fd15a5;
        exp_re_rom[398] = 'h7e2a2;
        exp_re_rom[399] = 'h46e6f;
        exp_re_rom[400] = 'h53f32;
        exp_re_rom[401] = 'hc2649;
        exp_re_rom[402] = 'h7f1c451;
        exp_re_rom[403] = 'h7fc29bb;
        exp_re_rom[404] = 'h7fe21a1;
        exp_re_rom[405] = 'h7ffb479;
        exp_re_rom[406] = 'h7fcd545;
        exp_re_rom[407] = 'h7fe6511;
        exp_re_rom[408] = 'h7feb2a5;
        exp_re_rom[409] = 'h7fe4b9d;
        exp_re_rom[410] = 'h192ac;
        exp_re_rom[411] = 'hc634;
        exp_re_rom[412] = 'h17c12;
        exp_re_rom[413] = 'h53262;
        exp_re_rom[414] = 'h7f506fd;
        exp_re_rom[415] = 'h7fbf4cf;
        exp_re_rom[416] = 'h7fca183;
        exp_re_rom[417] = 'h7fb12e1;
        exp_re_rom[418] = 'h45bd4;
        exp_re_rom[419] = 'h5aea;
        exp_re_rom[420] = 'h7ffcb0c;
        exp_re_rom[421] = 'h7ff7969;
        exp_re_rom[422] = 'hb0d;
        exp_re_rom[423] = 'h7ffa99c;
        exp_re_rom[424] = 'h7ff82b9;
        exp_re_rom[425] = 'h7ff14f9;
        exp_re_rom[426] = 'h12764;
        exp_re_rom[427] = 'h2451;
        exp_re_rom[428] = 'h1d1;
        exp_re_rom[429] = 'h7ffefa4;
        exp_re_rom[430] = 'h29e2;
        exp_re_rom[431] = 'h14d8;
        exp_re_rom[432] = 'h2145;
        exp_re_rom[433] = 'h4fe7;
        exp_re_rom[434] = 'h7ff85dc;
        exp_re_rom[435] = 'h96c;
        exp_re_rom[436] = 'h33f5;
        exp_re_rom[437] = 'h77f6;
        exp_re_rom[438] = 'h7ffbd0a;
        exp_re_rom[439] = 'h7045;
        exp_re_rom[440] = 'he6f7;
        exp_re_rom[441] = 'h23018;
        exp_re_rom[442] = 'h7fb7a8e;
        exp_re_rom[443] = 'h7ffe139;
        exp_re_rom[444] = 'h151af;
        exp_re_rom[445] = 'h52d6e;
        exp_re_rom[446] = 'h7ebe1f0;
        exp_re_rom[447] = 'h7fa956a;
        exp_re_rom[448] = 'h7fbd0a6;
        exp_re_rom[449] = 'h7fa9416;
        exp_re_rom[450] = 'h926bf;
        exp_re_rom[451] = 'hdee9;
        exp_re_rom[452] = 'h5305;
        exp_re_rom[453] = 'hf36e;
        exp_re_rom[454] = 'h7f9c986;
        exp_re_rom[455] = 'h7fe142b;
        exp_re_rom[456] = 'h7fe5a18;
        exp_re_rom[457] = 'h7fdfdc7;
        exp_re_rom[458] = 'h25d20;
        exp_re_rom[459] = 'h7ff9d80;
        exp_re_rom[460] = 'h7ff6597;
        exp_re_rom[461] = 'h7ff7257;
        exp_re_rom[462] = 'h7fdcf1c;
        exp_re_rom[463] = 'h7fec0f0;
        exp_re_rom[464] = 'h7feb7d6;
        exp_re_rom[465] = 'h7fe7f87;
        exp_re_rom[466] = 'h7ffcc33;
        exp_re_rom[467] = 'h7fe8f1f;
        exp_re_rom[468] = 'h7fe013c;
        exp_re_rom[469] = 'h7fc8068;
        exp_re_rom[470] = 'hbb32f;
        exp_re_rom[471] = 'h7542;
        exp_re_rom[472] = 'h7ff34cc;
        exp_re_rom[473] = 'h7fdc07f;
        exp_re_rom[474] = 'h92321;
        exp_re_rom[475] = 'h7ffb528;
        exp_re_rom[476] = 'h7fdd16e;
        exp_re_rom[477] = 'h7f94f33;
        exp_re_rom[478] = 'h36e17f;
        exp_re_rom[479] = 'h81df7;
        exp_re_rom[480] = 'h5d25e;
        exp_re_rom[481] = 'h6ee94;
        exp_re_rom[482] = 'h7e3fffd;
        exp_re_rom[483] = 'h7feff54;
        exp_re_rom[484] = 'h96d0;
        exp_re_rom[485] = 'h1fad7;
        exp_re_rom[486] = 'h7ef6764;
        exp_re_rom[487] = 'h7fecbc8;
        exp_re_rom[488] = 'h7ffa96d;
        exp_re_rom[489] = 'h3a48;
        exp_re_rom[490] = 'h7fa32b4;
        exp_re_rom[491] = 'h7ff818b;
        exp_re_rom[492] = 'h7ffd235;
        exp_re_rom[493] = 'h122e;
        exp_re_rom[494] = 'h7fc8cd3;
        exp_re_rom[495] = 'h7ffb936;
        exp_re_rom[496] = 'h7ffe0c3;
        exp_re_rom[497] = 'h7fff9d7;
        exp_re_rom[498] = 'h7ff0f2c;
        exp_re_rom[499] = 'h7fff801;
        exp_re_rom[500] = 'h965;
        exp_re_rom[501] = 'h1b6a;
        exp_re_rom[502] = 'h7fef231;
        exp_re_rom[503] = 'h1f85;
        exp_re_rom[504] = 'h3ca4;
        exp_re_rom[505] = 'h775e;
        exp_re_rom[506] = 'h7f0ce4d;
        exp_re_rom[507] = 'h7ffdae3;
        exp_re_rom[508] = 'h21ce;
        exp_re_rom[509] = 'h730e;
        exp_re_rom[510] = 'h7c6f835;
        exp_re_rom[511] = 'h7ffb0c3;
        exp_re_rom[512] = 'h7fffff6;
        exp_re_rom[513] = 'h3f11;
        exp_re_rom[514] = 'h1e93dc;
        exp_re_rom[515] = 'h7fffbbf;
        exp_re_rom[516] = 'h4317;
        exp_re_rom[517] = 'ha4db;
        exp_re_rom[518] = 'h175120;
        exp_re_rom[519] = 'h7ffd69b;
        exp_re_rom[520] = 'h61f9;
        exp_re_rom[521] = 'h12259;
        exp_re_rom[522] = 'h1f7ce1;
        exp_re_rom[523] = 'h7ff00f5;
        exp_re_rom[524] = 'h7fff583;
        exp_re_rom[525] = 'hef05;
        exp_re_rom[526] = 'h1af460;
        exp_re_rom[527] = 'h7fe5765;
        exp_re_rom[528] = 'h7ff761d;
        exp_re_rom[529] = 'h77d4;
        exp_re_rom[530] = 'h149323;
        exp_re_rom[531] = 'h7fdd719;
        exp_re_rom[532] = 'h7feefb8;
        exp_re_rom[533] = 'h7ffd2ba;
        exp_re_rom[534] = 'he4858;
        exp_re_rom[535] = 'h7fd571e;
        exp_re_rom[536] = 'h7fe2574;
        exp_re_rom[537] = 'h7fe6517;
        exp_re_rom[538] = 'h7fe5ffb;
        exp_re_rom[539] = 'h7fe94cd;
        exp_re_rom[540] = 'h7fe9538;
        exp_re_rom[541] = 'h7fe9de8;
        exp_re_rom[542] = 'hf352;
        exp_re_rom[543] = 'h7fd6401;
        exp_re_rom[544] = 'h7fcdd4b;
        exp_re_rom[545] = 'h7fae038;
        exp_re_rom[546] = 'h7da064d;
        exp_re_rom[547] = 'h4fa62;
        exp_re_rom[548] = 'h1ce37;
        exp_re_rom[549] = 'h8562;
        exp_re_rom[550] = 'h7fa644d;
        exp_re_rom[551] = 'h1e76d;
        exp_re_rom[552] = 'h12e4c;
        exp_re_rom[553] = 'h10920;
        exp_re_rom[554] = 'h2d0b6;
        exp_re_rom[555] = 'h7fffa8d;
        exp_re_rom[556] = 'h1fdf;
        exp_re_rom[557] = 'h1442;
        exp_re_rom[558] = 'h7ff5d63;
        exp_re_rom[559] = 'h5660;
        exp_re_rom[560] = 'h2d10;
        exp_re_rom[561] = 'h7fff9b0;
        exp_re_rom[562] = 'h7fde32e;
        exp_re_rom[563] = 'h10cd6;
        exp_re_rom[564] = 'hc955;
        exp_re_rom[565] = 'he236;
        exp_re_rom[566] = 'h2c379;
        exp_re_rom[567] = 'h7ffcf39;
        exp_re_rom[568] = 'h2098;
        exp_re_rom[569] = 'h12c8;
        exp_re_rom[570] = 'h7fdb8fa;
        exp_re_rom[571] = 'h21c20;
        exp_re_rom[572] = 'h2207f;
        exp_re_rom[573] = 'h3506e;
        exp_re_rom[574] = 'heeb30;
        exp_re_rom[575] = 'h7fc1e5d;
        exp_re_rom[576] = 'h7ff2582;
        exp_re_rom[577] = 'h10db6;
        exp_re_rom[578] = 'hcbfed;
        exp_re_rom[579] = 'h7f902ef;
        exp_re_rom[580] = 'h7fb76b4;
        exp_re_rom[581] = 'h7fac97c;
        exp_re_rom[582] = 'h7ee0e91;
        exp_re_rom[583] = 'h5a639;
        exp_re_rom[584] = 'h24e48;
        exp_re_rom[585] = 'h1e1fd;
        exp_re_rom[586] = 'h4e008;
        exp_re_rom[587] = 'h7fe9661;
        exp_re_rom[588] = 'h7ff72a8;
        exp_re_rom[589] = 'h7ff655e;
        exp_re_rom[590] = 'h7fcf931;
        exp_re_rom[591] = 'h22527;
        exp_re_rom[592] = 'h192d5;
        exp_re_rom[593] = 'h1fcac;
        exp_re_rom[594] = 'h59b57;
        exp_re_rom[595] = 'h7ff0526;
        exp_re_rom[596] = 'hd99c;
        exp_re_rom[597] = 'h277ec;
        exp_re_rom[598] = 'hb3ebf;
        exp_re_rom[599] = 'h7fa41eb;
        exp_re_rom[600] = 'h7fe0d57;
        exp_re_rom[601] = 'h7ff792d;
        exp_re_rom[602] = 'h2845a;
        exp_re_rom[603] = 'h7fe3c81;
        exp_re_rom[604] = 'h4ea4;
        exp_re_rom[605] = 'h2e349;
        exp_re_rom[606] = 'h11eae7;
        exp_re_rom[607] = 'h7f150c6;
        exp_re_rom[608] = 'h7f863cd;
        exp_re_rom[609] = 'h7f97ef7;
        exp_re_rom[610] = 'h7f6ce5a;
        exp_re_rom[611] = 'h7fe1acc;
        exp_re_rom[612] = 'h7fbd27a;
        exp_re_rom[613] = 'h7f97fe4;
        exp_re_rom[614] = 'h7ec7c82;
        exp_re_rom[615] = 'hb0991;
        exp_re_rom[616] = 'h39ba6;
        exp_re_rom[617] = 'h23f8e;
        exp_re_rom[618] = 'h3a4e7;
        exp_re_rom[619] = 'h7fdfa00;
        exp_re_rom[620] = 'h7ff0c12;
        exp_re_rom[621] = 'h7ff150c;
        exp_re_rom[622] = 'h7fe8eb2;
        exp_re_rom[623] = 'h7ffd942;
        exp_re_rom[624] = 'h7ff7010;
        exp_re_rom[625] = 'h7ff4994;
        exp_re_rom[626] = 'h7ff04b5;
        exp_re_rom[627] = 'h7ff7e6c;
        exp_re_rom[628] = 'h7ff4e81;
        exp_re_rom[629] = 'h7ff45bf;
        exp_re_rom[630] = 'h7ff8cff;
        exp_re_rom[631] = 'h7fe5e50;
        exp_re_rom[632] = 'h7fe7322;
        exp_re_rom[633] = 'h7fdf628;
        exp_re_rom[634] = 'h7fae6a7;
        exp_re_rom[635] = 'h449f4;
        exp_re_rom[636] = 'h1f986;
        exp_re_rom[637] = 'h2dfd6;
        exp_re_rom[638] = 'hb1eef;
        exp_re_rom[639] = 'h7f03467;
        exp_re_rom[640] = 'h7f7bfdb;
        exp_re_rom[641] = 'h7f74bee;
        exp_re_rom[642] = 'h7ee1573;
        exp_re_rom[643] = 'hbefcc;
        exp_re_rom[644] = 'h1563f;
        exp_re_rom[645] = 'h7fe07f7;
        exp_re_rom[646] = 'h7f6417a;
        exp_re_rom[647] = 'hc99d8;
        exp_re_rom[648] = 'h465ef;
        exp_re_rom[649] = 'h3061c;
        exp_re_rom[650] = 'h41b0c;
        exp_re_rom[651] = 'h7fcd834;
        exp_re_rom[652] = 'h7feaee7;
        exp_re_rom[653] = 'h7fe3518;
        exp_re_rom[654] = 'h7fafed0;
        exp_re_rom[655] = 'h638bb;
        exp_re_rom[656] = 'h1c068;
        exp_re_rom[657] = 'hc21c;
        exp_re_rom[658] = 'h7ffb440;
        exp_re_rom[659] = 'h1df11;
        exp_re_rom[660] = 'haea7;
        exp_re_rom[661] = 'h41ae;
        exp_re_rom[662] = 'h7ff83d6;
        exp_re_rom[663] = 'h17eaa;
        exp_re_rom[664] = 'h6cda;
        exp_re_rom[665] = 'h7fff974;
        exp_re_rom[666] = 'h7fec78c;
        exp_re_rom[667] = 'h3482e;
        exp_re_rom[668] = 'h16202;
        exp_re_rom[669] = 'h149bf;
        exp_re_rom[670] = 'h25960;
        exp_re_rom[671] = 'h7fccff1;
        exp_re_rom[672] = 'h7ff14d8;
        exp_re_rom[673] = 'h7ff41da;
        exp_re_rom[674] = 'h7fec2ea;
        exp_re_rom[675] = 'h179bb;
        exp_re_rom[676] = 'h3cee;
        exp_re_rom[677] = 'had4;
        exp_re_rom[678] = 'h7fff658;
        exp_re_rom[679] = 'h7ffd2ee;
        exp_re_rom[680] = 'h7ffcaf0;
        exp_re_rom[681] = 'h7ffb67c;
        exp_re_rom[682] = 'h7ff7cf1;
        exp_re_rom[683] = 'h6cb9;
        exp_re_rom[684] = 'h7ffe98c;
        exp_re_rom[685] = 'h7ffd172;
        exp_re_rom[686] = 'h7ffcb42;
        exp_re_rom[687] = 'h7ff8577;
        exp_re_rom[688] = 'h7ff9323;
        exp_re_rom[689] = 'h7ff846d;
        exp_re_rom[690] = 'h7ff5fbd;
        exp_re_rom[691] = 'h7ffe202;
        exp_re_rom[692] = 'h7ff8551;
        exp_re_rom[693] = 'h7ff66cd;
        exp_re_rom[694] = 'h7ff3d8d;
        exp_re_rom[695] = 'h7ff9bb3;
        exp_re_rom[696] = 'h7ff4124;
        exp_re_rom[697] = 'h7ff1d0e;
        exp_re_rom[698] = 'h7ff0ef6;
        exp_re_rom[699] = 'h7fdaf33;
        exp_re_rom[700] = 'h7fdc70c;
        exp_re_rom[701] = 'h7fcc931;
        exp_re_rom[702] = 'h7f9037e;
        exp_re_rom[703] = 'h128e08;
        exp_re_rom[704] = 'h33d4b;
        exp_re_rom[705] = 'h14e91;
        exp_re_rom[706] = 'h7fff783;
        exp_re_rom[707] = 'h40db9;
        exp_re_rom[708] = 'he7bb;
        exp_re_rom[709] = 'h2958;
        exp_re_rom[710] = 'h7fef27e;
        exp_re_rom[711] = 'h63590;
        exp_re_rom[712] = 'h1355d;
        exp_re_rom[713] = 'h4fb6;
        exp_re_rom[714] = 'h7febe07;
        exp_re_rom[715] = 'haf17a;
        exp_re_rom[716] = 'h319a1;
        exp_re_rom[717] = 'h2d904;
        exp_re_rom[718] = 'h496aa;
        exp_re_rom[719] = 'h7f0478a;
        exp_re_rom[720] = 'h7fda406;
        exp_re_rom[721] = 'h7fe9205;
        exp_re_rom[722] = 'h7fe7716;
        exp_re_rom[723] = 'h2f24c;
        exp_re_rom[724] = 'h7ffdfed;
        exp_re_rom[725] = 'h7ff8115;
        exp_re_rom[726] = 'h7fef40f;
        exp_re_rom[727] = 'h3c480;
        exp_re_rom[728] = 'h1216;
        exp_re_rom[729] = 'h7ff9816;
        exp_re_rom[730] = 'h7fefe06;
        exp_re_rom[731] = 'h374e0;
        exp_re_rom[732] = 'h7ff932b;
        exp_re_rom[733] = 'h7fea40f;
        exp_re_rom[734] = 'h7fc5549;
        exp_re_rom[735] = 'h1bfc6c;
        exp_re_rom[736] = 'h379f9;
        exp_re_rom[737] = 'h1ecb3;
        exp_re_rom[738] = 'h13cbd;
        exp_re_rom[739] = 'h34055;
        exp_re_rom[740] = 'h14439;
        exp_re_rom[741] = 'h1171c;
        exp_re_rom[742] = 'h11b6b;
        exp_re_rom[743] = 'h7fe6cd7;
        exp_re_rom[744] = 'h875b;
        exp_re_rom[745] = 'ha1dc;
        exp_re_rom[746] = 'hcc97;
        exp_re_rom[747] = 'h7fce0a2;
        exp_re_rom[748] = 'h3268;
        exp_re_rom[749] = 'h59a7;
        exp_re_rom[750] = 'h811f;
        exp_re_rom[751] = 'h7fd1214;
        exp_re_rom[752] = 'h1cdc;
        exp_re_rom[753] = 'h4095;
        exp_re_rom[754] = 'h6c31;
        exp_re_rom[755] = 'h7fb3c71;
        exp_re_rom[756] = 'h7fff831;
        exp_re_rom[757] = 'h2566;
        exp_re_rom[758] = 'h627e;
        exp_re_rom[759] = 'h7f4be0a;
        exp_re_rom[760] = 'h7ff98a5;
        exp_re_rom[761] = 'h7ffc75b;
        exp_re_rom[762] = 'h7ffd72b;
        exp_re_rom[763] = 'h7fe9360;
        exp_re_rom[764] = 'h7ffcadb;
        exp_re_rom[765] = 'h7ffc4d7;
        exp_re_rom[766] = 'h7ffaafb;
        exp_re_rom[767] = 'h2f5bd9;
        exp_re_rom[768] = 'h2;
        exp_re_rom[769] = 'h7ffde07;
        exp_re_rom[770] = 'h7ffc11a;
        exp_re_rom[771] = 'h7f6f942;
        exp_re_rom[772] = 'h7ffd49c;
        exp_re_rom[773] = 'h7ffa9aa;
        exp_re_rom[774] = 'h7ff5fc3;
        exp_re_rom[775] = 'h7eef70c;
        exp_re_rom[776] = 'h1c23;
        exp_re_rom[777] = 'h7ffad85;
        exp_re_rom[778] = 'h7ff18e1;
        exp_re_rom[779] = 'h7e990fc;
        exp_re_rom[780] = 'hc399;
        exp_re_rom[781] = 'h7fff86a;
        exp_re_rom[782] = 'h7fefc43;
        exp_re_rom[783] = 'h7e11dec;
        exp_re_rom[784] = 'h2c031;
        exp_re_rom[785] = 'h1e94d;
        exp_re_rom[786] = 'h22798;
        exp_re_rom[787] = 'h120201;
        exp_re_rom[788] = 'h7ff5f89;
        exp_re_rom[789] = 'h1e2b;
        exp_re_rom[790] = 'h8ef6;
        exp_re_rom[791] = 'h6566c;
        exp_re_rom[792] = 'h7ffa2ec;
        exp_re_rom[793] = 'h1812;
        exp_re_rom[794] = 'h843b;
        exp_re_rom[795] = 'h62461;
        exp_re_rom[796] = 'h7ff7a88;
        exp_re_rom[797] = 'h23a1;
        exp_re_rom[798] = 'h11109;
        exp_re_rom[799] = 'h100d37;
        exp_re_rom[800] = 'h7fcccd2;
        exp_re_rom[801] = 'h7fdd3d9;
        exp_re_rom[802] = 'h7fd9ab7;
        exp_re_rom[803] = 'h7f4925d;
        exp_re_rom[804] = 'hbfb2;
        exp_re_rom[805] = 'h7ffd792;
        exp_re_rom[806] = 'h7ff670e;
        exp_re_rom[807] = 'h7fc5f7b;
        exp_re_rom[808] = 'h4759;
        exp_re_rom[809] = 'h7ffe43a;
        exp_re_rom[810] = 'h7ffb88b;
        exp_re_rom[811] = 'h7ff2f01;
        exp_re_rom[812] = 'h7ffc2cd;
        exp_re_rom[813] = 'h7ffa4e6;
        exp_re_rom[814] = 'h7ff8f37;
        exp_re_rom[815] = 'h7ff454b;
        exp_re_rom[816] = 'h7ff8e0c;
        exp_re_rom[817] = 'h7ff76f4;
        exp_re_rom[818] = 'h7ff66c5;
        exp_re_rom[819] = 'h7ff8b81;
        exp_re_rom[820] = 'h7ff0abd;
        exp_re_rom[821] = 'h7fedac3;
        exp_re_rom[822] = 'h7fe524f;
        exp_re_rom[823] = 'h7f8fed7;
        exp_re_rom[824] = 'h13f41;
        exp_re_rom[825] = 'h59b8;
        exp_re_rom[826] = 'h8510;
        exp_re_rom[827] = 'h65240;
        exp_re_rom[828] = 'h7fbe295;
        exp_re_rom[829] = 'h7fc6386;
        exp_re_rom[830] = 'h7fae13b;
        exp_re_rom[831] = 'h7eb32dd;
        exp_re_rom[832] = 'h4fa4f;
        exp_re_rom[833] = 'heae4;
        exp_re_rom[834] = 'h7fecd0e;
        exp_re_rom[835] = 'h7f478eb;
        exp_re_rom[836] = 'h538fe;
        exp_re_rom[837] = 'h2a09e;
        exp_re_rom[838] = 'h242d7;
        exp_re_rom[839] = 'h60fb0;
        exp_re_rom[840] = 'h7fe03ae;
        exp_re_rom[841] = 'h7feddef;
        exp_re_rom[842] = 'h7feb22e;
        exp_re_rom[843] = 'h7fd09f6;
        exp_re_rom[844] = 'h7ff4a0a;
        exp_re_rom[845] = 'h7fe1601;
        exp_re_rom[846] = 'h7fc277e;
        exp_re_rom[847] = 'h7ef2403;
        exp_re_rom[848] = 'h74511;
        exp_re_rom[849] = 'h272d3;
        exp_re_rom[850] = 'h7787;
        exp_re_rom[851] = 'h7fa120e;
        exp_re_rom[852] = 'h55f83;
        exp_re_rom[853] = 'h312e2;
        exp_re_rom[854] = 'h2d515;
        exp_re_rom[855] = 'h62bce;
        exp_re_rom[856] = 'h7fe0609;
        exp_re_rom[857] = 'h7ff3c11;
        exp_re_rom[858] = 'h7ff168a;
        exp_re_rom[859] = 'h7fd3585;
        exp_re_rom[860] = 'h8c2c;
        exp_re_rom[861] = 'h7ff1c20;
        exp_re_rom[862] = 'h7fd57d5;
        exp_re_rom[863] = 'h7f35903;
        exp_re_rom[864] = 'h8d9e4;
        exp_re_rom[865] = 'h3cb6a;
        exp_re_rom[866] = 'h2662c;
        exp_re_rom[867] = 'h9aae;
        exp_re_rom[868] = 'h348b2;
        exp_re_rom[869] = 'h28a26;
        exp_re_rom[870] = 'h2abd5;
        exp_re_rom[871] = 'h54ae9;
        exp_re_rom[872] = 'h7fe69cc;
        exp_re_rom[873] = 'h7fff181;
        exp_re_rom[874] = 'h2196;
        exp_re_rom[875] = 'h7ffb302;
        exp_re_rom[876] = 'he64a;
        exp_re_rom[877] = 'h8394;
        exp_re_rom[878] = 'h4eb9;
        exp_re_rom[879] = 'h7ffc065;
        exp_re_rom[880] = 'hc508;
        exp_re_rom[881] = 'h4c18;
        exp_re_rom[882] = 'h7ffff30;
        exp_re_rom[883] = 'h7ff67f7;
        exp_re_rom[884] = 'h7ffd26c;
        exp_re_rom[885] = 'h7fed8cf;
        exp_re_rom[886] = 'h7fd0721;
        exp_re_rom[887] = 'h7f35fb0;
        exp_re_rom[888] = 'he733a;
        exp_re_rom[889] = 'h6bd94;
        exp_re_rom[890] = 'h63e03;
        exp_re_rom[891] = 'hc7576;
        exp_re_rom[892] = 'h7f6df3f;
        exp_re_rom[893] = 'h7fc57c4;
        exp_re_rom[894] = 'h7fb6c07;
        exp_re_rom[895] = 'h7f0e245;
        exp_re_rom[896] = 'h12b0c1;
        exp_re_rom[897] = 'h8279c;
        exp_re_rom[898] = 'h6bc43;
        exp_re_rom[899] = 'h86d73;
        exp_re_rom[900] = 'h1bcd6;
        exp_re_rom[901] = 'h4edbf;
        exp_re_rom[902] = 'h7d580;
        exp_re_rom[903] = 'h14a878;
        exp_re_rom[904] = 'h7eaf4b4;
        exp_re_rom[905] = 'h7f9db72;
        exp_re_rom[906] = 'h7fc8de8;
        exp_re_rom[907] = 'h7fd3cdd;
        exp_re_rom[908] = 'h7ff4dbc;
        exp_re_rom[909] = 'h7fef693;
        exp_re_rom[910] = 'h7feb156;
        exp_re_rom[911] = 'h7fca919;
        exp_re_rom[912] = 'h4f428;
        exp_re_rom[913] = 'h21c77;
        exp_re_rom[914] = 'h2019d;
        exp_re_rom[915] = 'h33051;
        exp_re_rom[916] = 'h7ff15bd;
        exp_re_rom[917] = 'h16937;
        exp_re_rom[918] = 'h32ad3;
        exp_re_rom[919] = 'ha241d;
        exp_re_rom[920] = 'h7ee656b;
        exp_re_rom[921] = 'h7f989ab;
        exp_re_rom[922] = 'h7fa890c;
        exp_re_rom[923] = 'h7f77312;
        exp_re_rom[924] = 'h6f926;
        exp_re_rom[925] = 'h1146;
        exp_re_rom[926] = 'h7fe08b5;
        exp_re_rom[927] = 'h7f8dad5;
        exp_re_rom[928] = 'he00ad;
        exp_re_rom[929] = 'h46e81;
        exp_re_rom[930] = 'h3182e;
        exp_re_rom[931] = 'h351da;
        exp_re_rom[932] = 'h7ff2af8;
        exp_re_rom[933] = 'hcc9d;
        exp_re_rom[934] = 'h1070b;
        exp_re_rom[935] = 'h17170;
        exp_re_rom[936] = 'h7ff65ed;
        exp_re_rom[937] = 'h5015;
        exp_re_rom[938] = 'h5604;
        exp_re_rom[939] = 'h7fff4d1;
        exp_re_rom[940] = 'h221ed;
        exp_re_rom[941] = 'h10d98;
        exp_re_rom[942] = 'he550;
        exp_re_rom[943] = 'hcc12;
        exp_re_rom[944] = 'hf9bf;
        exp_re_rom[945] = 'hd3bb;
        exp_re_rom[946] = 'hc032;
        exp_re_rom[947] = 'h85d8;
        exp_re_rom[948] = 'h1c1b7;
        exp_re_rom[949] = 'h10f34;
        exp_re_rom[950] = 'he7b0;
        exp_re_rom[951] = 'h94dd;
        exp_re_rom[952] = 'h24db5;
        exp_re_rom[953] = 'h135ee;
        exp_re_rom[954] = 'hc034;
        exp_re_rom[955] = 'h7fefb29;
        exp_re_rom[956] = 'hc7dcb;
        exp_re_rom[957] = 'h5ab42;
        exp_re_rom[958] = 'h6688a;
        exp_re_rom[959] = 'hc0e9e;
        exp_re_rom[960] = 'h7e2198e;
        exp_re_rom[961] = 'h7faf99c;
        exp_re_rom[962] = 'h7fd99e9;
        exp_re_rom[963] = 'h7fe26f9;
        exp_re_rom[964] = 'h313a7;
        exp_re_rom[965] = 'h103c0;
        exp_re_rom[966] = 'h176ea;
        exp_re_rom[967] = 'h34af7;
        exp_re_rom[968] = 'h7f51532;
        exp_re_rom[969] = 'h7fe494d;
        exp_re_rom[970] = 'h7ff3368;
        exp_re_rom[971] = 'h7ff42cc;
        exp_re_rom[972] = 'h39b05;
        exp_re_rom[973] = 'h17119;
        exp_re_rom[974] = 'h1ea66;
        exp_re_rom[975] = 'h3f02a;
        exp_re_rom[976] = 'h7f0f196;
        exp_re_rom[977] = 'h7fe1d5d;
        exp_re_rom[978] = 'h7ff764b;
        exp_re_rom[979] = 'h7db7;
        exp_re_rom[980] = 'h7fb5a50;
        exp_re_rom[981] = 'h7ff8a88;
        exp_re_rom[982] = 'h4921;
        exp_re_rom[983] = 'h1859a;
        exp_re_rom[984] = 'h7f5fbcc;
        exp_re_rom[985] = 'h7feb51b;
        exp_re_rom[986] = 'h7ff8f6d;
        exp_re_rom[987] = 'h4ac8;
        exp_re_rom[988] = 'h7fb8ffc;
        exp_re_rom[989] = 'h7ff9beb;
        exp_re_rom[990] = 'h4b51;
        exp_re_rom[991] = 'h19877;
        exp_re_rom[992] = 'h7f0d98e;
        exp_re_rom[993] = 'h7fe1286;
        exp_re_rom[994] = 'h7fefcd7;
        exp_re_rom[995] = 'h7ff9386;
        exp_re_rom[996] = 'h7fb6188;
        exp_re_rom[997] = 'h7ff0c3b;
        exp_re_rom[998] = 'h7ff5de6;
        exp_re_rom[999] = 'h7ffa6e0;
        exp_re_rom[1000] = 'h7fcbc71;
        exp_re_rom[1001] = 'h7ff4cf4;
        exp_re_rom[1002] = 'h7ff7b46;
        exp_re_rom[1003] = 'h7ff9dd3;
        exp_re_rom[1004] = 'h7fe6365;
        exp_re_rom[1005] = 'h7ff87c2;
        exp_re_rom[1006] = 'h7ff9ba5;
        exp_re_rom[1007] = 'h7ffa744;
        exp_re_rom[1008] = 'h7ffa8d5;
        exp_re_rom[1009] = 'h7ffb593;
        exp_re_rom[1010] = 'h7ffbad2;
        exp_re_rom[1011] = 'h7ffbc85;
        exp_re_rom[1012] = 'h5e1f;
        exp_re_rom[1013] = 'h7ffd34c;
        exp_re_rom[1014] = 'h7ffd2c3;
        exp_re_rom[1015] = 'h7ffd05f;
        exp_re_rom[1016] = 'h129c8;
        exp_re_rom[1017] = 'h7ffebee;
        exp_re_rom[1018] = 'h7ffea11;
        exp_re_rom[1019] = 'h7ffea39;
        exp_re_rom[1020] = 'hc598;
        exp_re_rom[1021] = 'h7fff70a;
        exp_re_rom[1022] = 'h7fff909;
        exp_re_rom[1023] = 'h7fffc4f;
    end
end
initial begin
    if (FFT_MODE) begin
        exp_im_rom[0] = 'h7fffeaa;
        exp_im_rom[1] = 'h7fffe52;
        exp_im_rom[2] = 'h7fffdcb;
        exp_im_rom[3] = 'h1a;
        exp_im_rom[4] = 'h1cd5d;
        exp_im_rom[5] = 'h7fff09b;
        exp_im_rom[6] = 'h7fff613;
        exp_im_rom[7] = 'h7ffff60;
        exp_im_rom[8] = 'h25b70;
        exp_im_rom[9] = 'h7ffd74d;
        exp_im_rom[10] = 'h7ffe1a6;
        exp_im_rom[11] = 'h7ffe77c;
        exp_im_rom[12] = 'h8ad0;
        exp_im_rom[13] = 'h7ffd752;
        exp_im_rom[14] = 'h7ffdac5;
        exp_im_rom[15] = 'h7ffdace;
        exp_im_rom[16] = 'h7ffd167;
        exp_im_rom[17] = 'h7ffd9cf;
        exp_im_rom[18] = 'h7ffd781;
        exp_im_rom[19] = 'h7ffd450;
        exp_im_rom[20] = 'h7ffc2f5;
        exp_im_rom[21] = 'h7ffcd4f;
        exp_im_rom[22] = 'h7ffc2c4;
        exp_im_rom[23] = 'h7ffa96e;
        exp_im_rom[24] = 'h7fdb2e7;
        exp_im_rom[25] = 'h7b4;
        exp_im_rom[26] = 'h7ffe0e4;
        exp_im_rom[27] = 'h7ffc4bf;
        exp_im_rom[28] = 'h7fedee5;
        exp_im_rom[29] = 'h7ffcd89;
        exp_im_rom[30] = 'h7ff89aa;
        exp_im_rom[31] = 'h7fee888;
        exp_im_rom[32] = 'h7f3cf42;
        exp_im_rom[33] = 'h248bc;
        exp_im_rom[34] = 'h1885b;
        exp_im_rom[35] = 'h1cbc5;
        exp_im_rom[36] = 'h9bdaa;
        exp_im_rom[37] = 'h7ff04a1;
        exp_im_rom[38] = 'h7ffdee5;
        exp_im_rom[39] = 'h4b0c;
        exp_im_rom[40] = 'h2d3c8;
        exp_im_rom[41] = 'h7ffb70f;
        exp_im_rom[42] = 'h3879;
        exp_im_rom[43] = 'hda69;
        exp_im_rom[44] = 'h78e7b;
        exp_im_rom[45] = 'h7fe26e3;
        exp_im_rom[46] = 'h7ff037c;
        exp_im_rom[47] = 'h7ff11b3;
        exp_im_rom[48] = 'h7fbaec5;
        exp_im_rom[49] = 'h15a32;
        exp_im_rom[50] = 'h1468b;
        exp_im_rom[51] = 'h242e6;
        exp_im_rom[52] = 'hde2fb;
        exp_im_rom[53] = 'h7fc5bf3;
        exp_im_rom[54] = 'h7fe7980;
        exp_im_rom[55] = 'h7ff53fd;
        exp_im_rom[56] = 'h1df1c;
        exp_im_rom[57] = 'h7fee851;
        exp_im_rom[58] = 'h7ffea6c;
        exp_im_rom[59] = 'h18179;
        exp_im_rom[60] = 'hfc7f9;
        exp_im_rom[61] = 'h7f88e24;
        exp_im_rom[62] = 'h7fb6194;
        exp_im_rom[63] = 'h7fba0d5;
        exp_im_rom[64] = 'h7f78e06;
        exp_im_rom[65] = 'h7fe81ff;
        exp_im_rom[66] = 'h7fce30d;
        exp_im_rom[67] = 'h7fab546;
        exp_im_rom[68] = 'h7e928fc;
        exp_im_rom[69] = 'h7a571;
        exp_im_rom[70] = 'h339d0;
        exp_im_rom[71] = 'h2a327;
        exp_im_rom[72] = 'h78985;
        exp_im_rom[73] = 'h7fd549c;
        exp_im_rom[74] = 'h7fea9a7;
        exp_im_rom[75] = 'h7fec748;
        exp_im_rom[76] = 'h7fdb7dc;
        exp_im_rom[77] = 'h7ffcf44;
        exp_im_rom[78] = 'h7ff6bbb;
        exp_im_rom[79] = 'h7ff46d7;
        exp_im_rom[80] = 'h7ff0986;
        exp_im_rom[81] = 'h7ff49d1;
        exp_im_rom[82] = 'h7ff2fc0;
        exp_im_rom[83] = 'h7ff2e65;
        exp_im_rom[84] = 'h7ffd46b;
        exp_im_rom[85] = 'h7fe1b22;
        exp_im_rom[86] = 'h7fe20fd;
        exp_im_rom[87] = 'h7fd95b7;
        exp_im_rom[88] = 'h7f9bdf5;
        exp_im_rom[89] = 'h18987;
        exp_im_rom[90] = 'h7ffdda4;
        exp_im_rom[91] = 'h7ff7fac;
        exp_im_rom[92] = 'h51be;
        exp_im_rom[93] = 'h7fd5804;
        exp_im_rom[94] = 'h7fd5569;
        exp_im_rom[95] = 'h7fc4963;
        exp_im_rom[96] = 'h7f5bc8e;
        exp_im_rom[97] = 'h3acfa;
        exp_im_rom[98] = 'h2e7;
        exp_im_rom[99] = 'h7fe6714;
        exp_im_rom[100] = 'h7f98da5;
        exp_im_rom[101] = 'h31253;
        exp_im_rom[102] = 'h213b;
        exp_im_rom[103] = 'h7fe996c;
        exp_im_rom[104] = 'h7f9568d;
        exp_im_rom[105] = 'h4c539;
        exp_im_rom[106] = 'h1af3d;
        exp_im_rom[107] = 'h12b87;
        exp_im_rom[108] = 'h34d7e;
        exp_im_rom[109] = 'h7fb9a0c;
        exp_im_rom[110] = 'h7fc7a88;
        exp_im_rom[111] = 'h7fadcd8;
        exp_im_rom[112] = 'h7f0bbc5;
        exp_im_rom[113] = 'ha70ec;
        exp_im_rom[114] = 'h2d503;
        exp_im_rom[115] = 'h84e5;
        exp_im_rom[116] = 'h7fc52a6;
        exp_im_rom[117] = 'h4b69e;
        exp_im_rom[118] = 'h17c70;
        exp_im_rom[119] = 'h7fffe1a;
        exp_im_rom[120] = 'h7fbad24;
        exp_im_rom[121] = 'h6a17b;
        exp_im_rom[122] = 'h36738;
        exp_im_rom[123] = 'h3aaf2;
        exp_im_rom[124] = 'ha6452;
        exp_im_rom[125] = 'h7f2e360;
        exp_im_rom[126] = 'h7f838f1;
        exp_im_rom[127] = 'h7f5ab82;
        exp_im_rom[128] = 'h7e2cc71;
        exp_im_rom[129] = 'h1d920d;
        exp_im_rom[130] = 'ha1290;
        exp_im_rom[131] = 'h61199;
        exp_im_rom[132] = 'h31755;
        exp_im_rom[133] = 'h7688c;
        exp_im_rom[134] = 'h5b18d;
        exp_im_rom[135] = 'h64875;
        exp_im_rom[136] = 'hc306a;
        exp_im_rom[137] = 'h7f6dde1;
        exp_im_rom[138] = 'h7fe24e3;
        exp_im_rom[139] = 'h7ff23e9;
        exp_im_rom[140] = 'h7fe5dc6;
        exp_im_rom[141] = 'h2d516;
        exp_im_rom[142] = 'h154ee;
        exp_im_rom[143] = 'h11702;
        exp_im_rom[144] = 'hfc45;
        exp_im_rom[145] = 'hf0ac;
        exp_im_rom[146] = 'hdfc3;
        exp_im_rom[147] = 'hcc37;
        exp_im_rom[148] = 'h97d4;
        exp_im_rom[149] = 'h12422;
        exp_im_rom[150] = 'hcb5f;
        exp_im_rom[151] = 'h84cc;
        exp_im_rom[152] = 'h7ff63a5;
        exp_im_rom[153] = 'h416d7;
        exp_im_rom[154] = 'h2486f;
        exp_im_rom[155] = 'h24883;
        exp_im_rom[156] = 'h36809;
        exp_im_rom[157] = 'h7feab92;
        exp_im_rom[158] = 'h10ffa;
        exp_im_rom[159] = 'h21aee;
        exp_im_rom[160] = 'h55ff6;
        exp_im_rom[161] = 'h7f77484;
        exp_im_rom[162] = 'h7fdc793;
        exp_im_rom[163] = 'h7fea113;
        exp_im_rom[164] = 'h7fe48c8;
        exp_im_rom[165] = 'h26d19;
        exp_im_rom[166] = 'h103bd;
        exp_im_rom[167] = 'h176b1;
        exp_im_rom[168] = 'h43f0d;
        exp_im_rom[169] = 'h7f595ac;
        exp_im_rom[170] = 'h7fc5807;
        exp_im_rom[171] = 'h7fcb538;
        exp_im_rom[172] = 'h7fab1f5;
        exp_im_rom[173] = 'h69a44;
        exp_im_rom[174] = 'h6665;
        exp_im_rom[175] = 'h7ff03bd;
        exp_im_rom[176] = 'h7fc608a;
        exp_im_rom[177] = 'h8c7e5;
        exp_im_rom[178] = 'h1eec8;
        exp_im_rom[179] = 'hc0a9;
        exp_im_rom[180] = 'h7ff93a1;
        exp_im_rom[181] = 'h366d4;
        exp_im_rom[182] = 'hd2fb;
        exp_im_rom[183] = 'h18c2;
        exp_im_rom[184] = 'h7fed303;
        exp_im_rom[185] = 'h4591f;
        exp_im_rom[186] = 'h8722;
        exp_im_rom[187] = 'h7ff1475;
        exp_im_rom[188] = 'h7fb014c;
        exp_im_rom[189] = 'h1584ca;
        exp_im_rom[190] = 'h65030;
        exp_im_rom[191] = 'h51d70;
        exp_im_rom[192] = 'h6b17b;
        exp_im_rom[193] = 'h7f62d37;
        exp_im_rom[194] = 'h7ffc457;
        exp_im_rom[195] = 'hd2c2;
        exp_im_rom[196] = 'h19e08;
        exp_im_rom[197] = 'h7fe2eeb;
        exp_im_rom[198] = 'h95e3;
        exp_im_rom[199] = 'h10663;
        exp_im_rom[200] = 'h1afa2;
        exp_im_rom[201] = 'h7fd9f62;
        exp_im_rom[202] = 'h7f4c;
        exp_im_rom[203] = 'h1114e;
        exp_im_rom[204] = 'h22d4d;
        exp_im_rom[205] = 'h7f95b88;
        exp_im_rom[206] = 'h7ff59ad;
        exp_im_rom[207] = 'h7fff785;
        exp_im_rom[208] = 'h59fb;
        exp_im_rom[209] = 'h7ff01d7;
        exp_im_rom[210] = 'h261c;
        exp_im_rom[211] = 'h6205;
        exp_im_rom[212] = 'hcb3f;
        exp_im_rom[213] = 'h7fd05ff;
        exp_im_rom[214] = 'h7ffbe84;
        exp_im_rom[215] = 'h7fff2e6;
        exp_im_rom[216] = 'h7fff7c8;
        exp_im_rom[217] = 'ha975;
        exp_im_rom[218] = 'h2150;
        exp_im_rom[219] = 'h7fff37a;
        exp_im_rom[220] = 'h7ff5210;
        exp_im_rom[221] = 'h8c003;
        exp_im_rom[222] = 'h1c9f1;
        exp_im_rom[223] = 'h1941f;
        exp_im_rom[224] = 'h228fd;
        exp_im_rom[225] = 'h7f70f75;
        exp_im_rom[226] = 'h7ffb92f;
        exp_im_rom[227] = 'h4860;
        exp_im_rom[228] = 'hb3e6;
        exp_im_rom[229] = 'h7fc9c32;
        exp_im_rom[230] = 'h1e35;
        exp_im_rom[231] = 'h6e34;
        exp_im_rom[232] = 'hd6ef;
        exp_im_rom[233] = 'h7fa79cd;
        exp_im_rom[234] = 'h7ffece8;
        exp_im_rom[235] = 'h3f61;
        exp_im_rom[236] = 'h7cb6;
        exp_im_rom[237] = 'h7fe9898;
        exp_im_rom[238] = 'h8df2;
        exp_im_rom[239] = 'hfa68;
        exp_im_rom[240] = 'h21395;
        exp_im_rom[241] = 'h7df394f;
        exp_im_rom[242] = 'h7fe41c6;
        exp_im_rom[243] = 'h7ff2fcb;
        exp_im_rom[244] = 'h7ffa080;
        exp_im_rom[245] = 'h7f92159;
        exp_im_rom[246] = 'h7ff426a;
        exp_im_rom[247] = 'h7ff5c01;
        exp_im_rom[248] = 'h7ff2cad;
        exp_im_rom[249] = 'h1213ff;
        exp_im_rom[250] = 'h3a7d;
        exp_im_rom[251] = 'h7fff3b8;
        exp_im_rom[252] = 'h7ffb42f;
        exp_im_rom[253] = 'h1e9de8;
        exp_im_rom[254] = 'h5d27;
        exp_im_rom[255] = 'h2658;
        exp_im_rom[256] = 'h10;
        exp_im_rom[257] = 'h7d74a32;
        exp_im_rom[258] = 'h3b1d;
        exp_im_rom[259] = 'h15f3;
        exp_im_rom[260] = 'h7ffe4e2;
        exp_im_rom[261] = 'h7f01077;
        exp_im_rom[262] = 'h7951;
        exp_im_rom[263] = 'h45a5;
        exp_im_rom[264] = 'h1e32;
        exp_im_rom[265] = 'h7fa82e8;
        exp_im_rom[266] = 'h7a7b;
        exp_im_rom[267] = 'h5bc5;
        exp_im_rom[268] = 'h5056;
        exp_im_rom[269] = 'h5494;
        exp_im_rom[270] = 'h416a;
        exp_im_rom[271] = 'h3898;
        exp_im_rom[272] = 'h1ff7;
        exp_im_rom[273] = 'h7fcffc7;
        exp_im_rom[274] = 'h9aa8;
        exp_im_rom[275] = 'h83ef;
        exp_im_rom[276] = 'h8d55;
        exp_im_rom[277] = 'h1cbd4;
        exp_im_rom[278] = 'h6c51;
        exp_im_rom[279] = 'ha125;
        exp_im_rom[280] = 'h112a9;
        exp_im_rom[281] = 'ha237d;
        exp_im_rom[282] = 'h7ff289d;
        exp_im_rom[283] = 'h7ffcc7f;
        exp_im_rom[284] = 'h343d;
        exp_im_rom[285] = 'h4eab2;
        exp_im_rom[286] = 'h7ff1422;
        exp_im_rom[287] = 'h7ff671b;
        exp_im_rom[288] = 'h7ff64f1;
        exp_im_rom[289] = 'h7fd8e37;
        exp_im_rom[290] = 'h7fffc01;
        exp_im_rom[291] = 'h7ffc54c;
        exp_im_rom[292] = 'h7ff9207;
        exp_im_rom[293] = 'h7fd73a1;
        exp_im_rom[294] = 'h29c5;
        exp_im_rom[295] = 'h7ffd974;
        exp_im_rom[296] = 'h7ff8f77;
        exp_im_rom[297] = 'h7fcec00;
        exp_im_rom[298] = 'h62da;
        exp_im_rom[299] = 'h7fff6b1;
        exp_im_rom[300] = 'h7ffa61a;
        exp_im_rom[301] = 'h7fd8e91;
        exp_im_rom[302] = 'h36f0;
        exp_im_rom[303] = 'h7ffb7b4;
        exp_im_rom[304] = 'h7ff2297;
        exp_im_rom[305] = 'h7fa2827;
        exp_im_rom[306] = 'h11ba6;
        exp_im_rom[307] = 'ha84;
        exp_im_rom[308] = 'h7ff0d51;
        exp_im_rom[309] = 'h7f6f0dc;
        exp_im_rom[310] = 'h31556;
        exp_im_rom[311] = 'h1af51;
        exp_im_rom[312] = 'h18314;
        exp_im_rom[313] = 'h4d9d0;
        exp_im_rom[314] = 'h7fe90cc;
        exp_im_rom[315] = 'h7fea961;
        exp_im_rom[316] = 'h7fd5178;
        exp_im_rom[317] = 'h7ef2d66;
        exp_im_rom[318] = 'h6740b;
        exp_im_rom[319] = 'h36b74;
        exp_im_rom[320] = 'h2cb6b;
        exp_im_rom[321] = 'h42552;
        exp_im_rom[322] = 'h133ab;
        exp_im_rom[323] = 'h1b3d5;
        exp_im_rom[324] = 'h25885;
        exp_im_rom[325] = 'h7d695;
        exp_im_rom[326] = 'h7fe1831;
        exp_im_rom[327] = 'h7ff8083;
        exp_im_rom[328] = 'h7ffb4cb;
        exp_im_rom[329] = 'h7fe9ecd;
        exp_im_rom[330] = 'hdcba;
        exp_im_rom[331] = 'h777e;
        exp_im_rom[332] = 'h3722;
        exp_im_rom[333] = 'h7fedf15;
        exp_im_rom[334] = 'h13bd8;
        exp_im_rom[335] = 'hba93;
        exp_im_rom[336] = 'h7859;
        exp_im_rom[337] = 'h7ffaca9;
        exp_im_rom[338] = 'hbe2c;
        exp_im_rom[339] = 'h2841;
        exp_im_rom[340] = 'h7ff3198;
        exp_im_rom[341] = 'h7f884fa;
        exp_im_rom[342] = 'h61ccc;
        exp_im_rom[343] = 'h3a823;
        exp_im_rom[344] = 'h39488;
        exp_im_rom[345] = 'h7557f;
        exp_im_rom[346] = 'h7fe9dda;
        exp_im_rom[347] = 'h190e;
        exp_im_rom[348] = 'h7ffcdbf;
        exp_im_rom[349] = 'h7faa8e8;
        exp_im_rom[350] = 'h72492;
        exp_im_rom[351] = 'h548cc;
        exp_im_rom[352] = 'h673e3;
        exp_im_rom[353] = 'h10bf1b;
        exp_im_rom[354] = 'h7f9beea;
        exp_im_rom[355] = 'h7ff9774;
        exp_im_rom[356] = 'h203c3;
        exp_im_rom[357] = 'h99db4;
        exp_im_rom[358] = 'h7f9cce1;
        exp_im_rom[359] = 'h7fe28a7;
        exp_im_rom[360] = 'h7ff9c1f;
        exp_im_rom[361] = 'h24cd7;
        exp_im_rom[362] = 'h7fd9160;
        exp_im_rom[363] = 'h7ff456e;
        exp_im_rom[364] = 'h2932;
        exp_im_rom[365] = 'h312ca;
        exp_im_rom[366] = 'h7fc58b2;
        exp_im_rom[367] = 'h7fe24c4;
        exp_im_rom[368] = 'h7fe41d5;
        exp_im_rom[369] = 'h7fc88b2;
        exp_im_rom[370] = 'h16f07;
        exp_im_rom[371] = 'h7ffc810;
        exp_im_rom[372] = 'h7fe825f;
        exp_im_rom[373] = 'h7f7dd30;
        exp_im_rom[374] = 'hb0839;
        exp_im_rom[375] = 'h66fc5;
        exp_im_rom[376] = 'h78660;
        exp_im_rom[377] = 'h12eea2;
        exp_im_rom[378] = 'h7f0f310;
        exp_im_rom[379] = 'h7faf527;
        exp_im_rom[380] = 'h7fc41e7;
        exp_im_rom[381] = 'h7f89ab7;
        exp_im_rom[382] = 'h763f1;
        exp_im_rom[383] = 'h3d7c2;
        exp_im_rom[384] = 'h4ac7d;
        exp_im_rom[385] = 'hbde92;
        exp_im_rom[386] = 'h7f58c8d;
        exp_im_rom[387] = 'h7fd6524;
        exp_im_rom[388] = 'h7ffa777;
        exp_im_rom[389] = 'h444b4;
        exp_im_rom[390] = 'h7f79251;
        exp_im_rom[391] = 'h7fc24f6;
        exp_im_rom[392] = 'h7fcb3b4;
        exp_im_rom[393] = 'h7faf729;
        exp_im_rom[394] = 'h295aa;
        exp_im_rom[395] = 'hc40;
        exp_im_rom[396] = 'h7ff99a0;
        exp_im_rom[397] = 'h7ff1db0;
        exp_im_rom[398] = 'h57e4;
        exp_im_rom[399] = 'h7ffcd47;
        exp_im_rom[400] = 'h7ff99d2;
        exp_im_rom[401] = 'h7ff0518;
        exp_im_rom[402] = 'h108af;
        exp_im_rom[403] = 'h3748;
        exp_im_rom[404] = 'h85d;
        exp_im_rom[405] = 'h7ffbfaa;
        exp_im_rom[406] = 'ha634;
        exp_im_rom[407] = 'h469e;
        exp_im_rom[408] = 'h410a;
        exp_im_rom[409] = 'h88b9;
        exp_im_rom[410] = 'h7fee651;
        exp_im_rom[411] = 'h7ff4a42;
        exp_im_rom[412] = 'h7fec681;
        exp_im_rom[413] = 'h7fbed43;
        exp_im_rom[414] = 'h8ccd9;
        exp_im_rom[415] = 'h379a4;
        exp_im_rom[416] = 'h331d6;
        exp_im_rom[417] = 'h54709;
        exp_im_rom[418] = 'h7fa8c8a;
        exp_im_rom[419] = 'h7ff66a5;
        exp_im_rom[420] = 'h3600;
        exp_im_rom[421] = 'hcd8a;
        exp_im_rom[422] = 'h7ffdfa7;
        exp_im_rom[423] = 'hb38e;
        exp_im_rom[424] = 'h135de;
        exp_im_rom[425] = 'h2a552;
        exp_im_rom[426] = 'h7fc57e1;
        exp_im_rom[427] = 'h7ffac32;
        exp_im_rom[428] = 'h56ad;
        exp_im_rom[429] = 'h107aa;
        exp_im_rom[430] = 'h7ff6159;
        exp_im_rom[431] = 'hb738;
        exp_im_rom[432] = 'h17078;
        exp_im_rom[433] = 'h36e32;
        exp_im_rom[434] = 'h7f98fd8;
        exp_im_rom[435] = 'h7ff18a1;
        exp_im_rom[436] = 'h1793;
        exp_im_rom[437] = 'h1135f;
        exp_im_rom[438] = 'h7fe6f41;
        exp_im_rom[439] = 'h9648;
        exp_im_rom[440] = 'h196c6;
        exp_im_rom[441] = 'h41351;
        exp_im_rom[442] = 'h7f70565;
        exp_im_rom[443] = 'h7ff4e01;
        exp_im_rom[444] = 'h18055;
        exp_im_rom[445] = 'h686d7;
        exp_im_rom[446] = 'h7e70c4c;
        exp_im_rom[447] = 'h7f99974;
        exp_im_rom[448] = 'h7fb66ee;
        exp_im_rom[449] = 'h7faaf0d;
        exp_im_rom[450] = 'h71e0b;
        exp_im_rom[451] = 'h42e8;
        exp_im_rom[452] = 'h7ffd6f8;
        exp_im_rom[453] = 'h331a;
        exp_im_rom[454] = 'h7fc50a0;
        exp_im_rom[455] = 'h7febb85;
        exp_im_rom[456] = 'h7fef6b3;
        exp_im_rom[457] = 'h7feeea6;
        exp_im_rom[458] = 'h5f2f;
        exp_im_rom[459] = 'h7ff8fe1;
        exp_im_rom[460] = 'h7ff8a9b;
        exp_im_rom[461] = 'h7ff9506;
        exp_im_rom[462] = 'h7ff7372;
        exp_im_rom[463] = 'h7ff9b74;
        exp_im_rom[464] = 'h7ffab97;
        exp_im_rom[465] = 'h7ffbecf;
        exp_im_rom[466] = 'h7ffb146;
        exp_im_rom[467] = 'h7ffe317;
        exp_im_rom[468] = 'h1206;
        exp_im_rom[469] = 'h8cb6;
        exp_im_rom[470] = 'h7fc1fa9;
        exp_im_rom[471] = 'h7ff8210;
        exp_im_rom[472] = 'h7ffffe8;
        exp_im_rom[473] = 'hbb73;
        exp_im_rom[474] = 'h7fac85e;
        exp_im_rom[475] = 'h7ffd6d5;
        exp_im_rom[476] = 'h11e49;
        exp_im_rom[477] = 'h49e45;
        exp_im_rom[478] = 'h7d29c9a;
        exp_im_rom[479] = 'h7f849d7;
        exp_im_rom[480] = 'h7f9d10f;
        exp_im_rom[481] = 'h7f7fb47;
        exp_im_rom[482] = 'h21bd1a;
        exp_im_rom[483] = 'hf5d8;
        exp_im_rom[484] = 'h7feb688;
        exp_im_rom[485] = 'h7fc4652;
        exp_im_rom[486] = 'h1e9b60;
        exp_im_rom[487] = 'h21399;
        exp_im_rom[488] = 'h508d;
        exp_im_rom[489] = 'h7fed1f5;
        exp_im_rom[490] = 'h12863b;
        exp_im_rom[491] = 'h149b4;
        exp_im_rom[492] = 'h1807;
        exp_im_rom[493] = 'h7fe82f4;
        exp_im_rom[494] = 'h2199ca;
        exp_im_rom[495] = 'h2f4e7;
        exp_im_rom[496] = 'h1f046;
        exp_im_rom[497] = 'h1d162;
        exp_im_rom[498] = 'h7f78399;
        exp_im_rom[499] = 'h71d6;
        exp_im_rom[500] = 'ha252;
        exp_im_rom[501] = 'hc0fe;
        exp_im_rom[502] = 'h7fcc558;
        exp_im_rom[503] = 'h8813;
        exp_im_rom[504] = 'hb742;
        exp_im_rom[505] = 'h118f3;
        exp_im_rom[506] = 'h7e3a889;
        exp_im_rom[507] = 'h7ffd248;
        exp_im_rom[508] = 'h3e5c;
        exp_im_rom[509] = 'ha34e;
        exp_im_rom[510] = 'h7ba870b;
        exp_im_rom[511] = 'h7ffaaee;
        exp_im_rom[512] = 'h6;
        exp_im_rom[513] = 'h3742;
        exp_im_rom[514] = 'h19149d;
        exp_im_rom[515] = 'h7fff7d2;
        exp_im_rom[516] = 'h268f;
        exp_im_rom[517] = 'h5b71;
        exp_im_rom[518] = 'hc6e2d;
        exp_im_rom[519] = 'h7ffe350;
        exp_im_rom[520] = 'h1ecc;
        exp_im_rom[521] = 'h5d8b;
        exp_im_rom[522] = 'h9827c;
        exp_im_rom[523] = 'h7ffb4f0;
        exp_im_rom[524] = 'h7fff274;
        exp_im_rom[525] = 'h17d4;
        exp_im_rom[526] = 'h29bf3;
        exp_im_rom[527] = 'h7ffdf6a;
        exp_im_rom[528] = 'h7fff447;
        exp_im_rom[529] = 'h7ffee95;
        exp_im_rom[530] = 'h7fdede3;
        exp_im_rom[531] = 'h46fc;
        exp_im_rom[532] = 'h2b83;
        exp_im_rom[533] = 'h143;
        exp_im_rom[534] = 'h7fba166;
        exp_im_rom[535] = 'heae6;
        exp_im_rom[536] = 'hbcad;
        exp_im_rom[537] = 'hbb6a;
        exp_im_rom[538] = 'hd89e;
        exp_im_rom[539] = 'hd551;
        exp_im_rom[540] = 'hef8d;
        exp_im_rom[541] = 'h10583;
        exp_im_rom[542] = 'h7ff3956;
        exp_im_rom[543] = 'h260be;
        exp_im_rom[544] = 'h328c0;
        exp_im_rom[545] = 'h5b0a8;
        exp_im_rom[546] = 'h2e52d5;
        exp_im_rom[547] = 'h7f95af7;
        exp_im_rom[548] = 'h7fd62c6;
        exp_im_rom[549] = 'h7ff3e7d;
        exp_im_rom[550] = 'haa26b;
        exp_im_rom[551] = 'h7fc275a;
        exp_im_rom[552] = 'h7fd6036;
        exp_im_rom[553] = 'h7fd64dd;
        exp_im_rom[554] = 'h7f71707;
        exp_im_rom[555] = 'h924f;
        exp_im_rom[556] = 'h991;
        exp_im_rom[557] = 'h6cfb;
        exp_im_rom[558] = 'h8014e;
        exp_im_rom[559] = 'h7fc7a41;
        exp_im_rom[560] = 'h7fcffa7;
        exp_im_rom[561] = 'h7fbaa24;
        exp_im_rom[562] = 'h7e88125;
        exp_im_rom[563] = 'h5a0ba;
        exp_im_rom[564] = 'h2cc1f;
        exp_im_rom[565] = 'h28c51;
        exp_im_rom[566] = 'h83f16;
        exp_im_rom[567] = 'h7feaf2d;
        exp_im_rom[568] = 'h7ff9578;
        exp_im_rom[569] = 'h7ff7a21;
        exp_im_rom[570] = 'h7fb18cc;
        exp_im_rom[571] = 'h2e7c7;
        exp_im_rom[572] = 'h29757;
        exp_im_rom[573] = 'h3e526;
        exp_im_rom[574] = 'h119ea0;
        exp_im_rom[575] = 'h7fb2b97;
        exp_im_rom[576] = 'h7fe9be4;
        exp_im_rom[577] = 'h6cc7;
        exp_im_rom[578] = 'h9f077;
        exp_im_rom[579] = 'h7fa4c18;
        exp_im_rom[580] = 'h7fc73d2;
        exp_im_rom[581] = 'h7fc5c63;
        exp_im_rom[582] = 'h7f5e530;
        exp_im_rom[583] = 'h22877;
        exp_im_rom[584] = 'h70ab;
        exp_im_rom[585] = 'h2828;
        exp_im_rom[586] = 'hf58f;
        exp_im_rom[587] = 'h7ff1f76;
        exp_im_rom[588] = 'h7ff5cb6;
        exp_im_rom[589] = 'h7ff608c;
        exp_im_rom[590] = 'h7ff2993;
        exp_im_rom[591] = 'h7ff8f13;
        exp_im_rom[592] = 'h7ff7216;
        exp_im_rom[593] = 'h7ff56d7;
        exp_im_rom[594] = 'h7fedff4;
        exp_im_rom[595] = 'h7ff8fab;
        exp_im_rom[596] = 'h7ff3c29;
        exp_im_rom[597] = 'h7fec5c4;
        exp_im_rom[598] = 'h7fbf71d;
        exp_im_rom[599] = 'h16a4f;
        exp_im_rom[600] = 'h2645;
        exp_im_rom[601] = 'h7ff9291;
        exp_im_rom[602] = 'h7fdf4d2;
        exp_im_rom[603] = 'h55d6;
        exp_im_rom[604] = 'h7ff0bf2;
        exp_im_rom[605] = 'h7fd14ac;
        exp_im_rom[606] = 'h7f07c47;
        exp_im_rom[607] = 'hc764b;
        exp_im_rom[608] = 'h6b8b0;
        exp_im_rom[609] = 'h63d84;
        exp_im_rom[610] = 'ha3661;
        exp_im_rom[611] = 'h180a6;
        exp_im_rom[612] = 'h52061;
        exp_im_rom[613] = 'h9a1c1;
        exp_im_rom[614] = 'h2330a1;
        exp_im_rom[615] = 'h7e737fe;
        exp_im_rom[616] = 'h7f5af87;
        exp_im_rom[617] = 'h7f7e867;
        exp_im_rom[618] = 'h7f1e7fb;
        exp_im_rom[619] = 'h59d69;
        exp_im_rom[620] = 'h1c0d4;
        exp_im_rom[621] = 'h23256;
        exp_im_rom[622] = 'h8be30;
        exp_im_rom[623] = 'h7f774e2;
        exp_im_rom[624] = 'h7fc0655;
        exp_im_rom[625] = 'h7fcc4fa;
        exp_im_rom[626] = 'h7fb9527;
        exp_im_rom[627] = 'h3993;
        exp_im_rom[628] = 'h7ff3274;
        exp_im_rom[629] = 'h7ff3470;
        exp_im_rom[630] = 'h3e6c;
        exp_im_rom[631] = 'h7fce40c;
        exp_im_rom[632] = 'h7fd80a0;
        exp_im_rom[633] = 'h7fcc631;
        exp_im_rom[634] = 'h7f76a4e;
        exp_im_rom[635] = 'h80116;
        exp_im_rom[636] = 'h3b714;
        exp_im_rom[637] = 'h48f38;
        exp_im_rom[638] = 'he2b6f;
        exp_im_rom[639] = 'h7ef225a;
        exp_im_rom[640] = 'h7f842b1;
        exp_im_rom[641] = 'h7f893e3;
        exp_im_rom[642] = 'h7f1b8d0;
        exp_im_rom[643] = 'h93dd9;
        exp_im_rom[644] = 'h13f9b;
        exp_im_rom[645] = 'h7ff24d0;
        exp_im_rom[646] = 'h7fb1641;
        exp_im_rom[647] = 'h63a7f;
        exp_im_rom[648] = 'h210ae;
        exp_im_rom[649] = 'h14d2b;
        exp_im_rom[650] = 'h17151;
        exp_im_rom[651] = 'h7ff6287;
        exp_im_rom[652] = 'h7ffe480;
        exp_im_rom[653] = 'h7ffde58;
        exp_im_rom[654] = 'h7ff9f2e;
        exp_im_rom[655] = 'h66bc;
        exp_im_rom[656] = 'h1397;
        exp_im_rom[657] = 'h53a;
        exp_im_rom[658] = 'h1173;
        exp_im_rom[659] = 'h7ffbe19;
        exp_im_rom[660] = 'h7ffdd90;
        exp_im_rom[661] = 'h7ffeafc;
        exp_im_rom[662] = 'h1bff;
        exp_im_rom[663] = 'h7ff6846;
        exp_im_rom[664] = 'h7ffbebd;
        exp_im_rom[665] = 'h7ffe94d;
        exp_im_rom[666] = 'h8745;
        exp_im_rom[667] = 'h7fde285;
        exp_im_rom[668] = 'h7fee6dd;
        exp_im_rom[669] = 'h7fed7c8;
        exp_im_rom[670] = 'h7fdd71a;
        exp_im_rom[671] = 'h29fd2;
        exp_im_rom[672] = 'h9e22;
        exp_im_rom[673] = 'h7a7e;
        exp_im_rom[674] = 'h11f75;
        exp_im_rom[675] = 'h7fd92bd;
        exp_im_rom[676] = 'h7ff25a8;
        exp_im_rom[677] = 'h7ff5d1d;
        exp_im_rom[678] = 'h7ff6c55;
        exp_im_rom[679] = 'h7ffa02b;
        exp_im_rom[680] = 'h7ffa14b;
        exp_im_rom[681] = 'h7ffc65a;
        exp_im_rom[682] = 'h7399;
        exp_im_rom[683] = 'h7fcc6d6;
        exp_im_rom[684] = 'h7fe7a5d;
        exp_im_rom[685] = 'h7fe893e;
        exp_im_rom[686] = 'h7fdf4e7;
        exp_im_rom[687] = 'h14789;
        exp_im_rom[688] = 'h7ff77fc;
        exp_im_rom[689] = 'h7ff07ab;
        exp_im_rom[690] = 'h7fe2a5c;
        exp_im_rom[691] = 'h2499b;
        exp_im_rom[692] = 'h7fff183;
        exp_im_rom[693] = 'h7ff876e;
        exp_im_rom[694] = 'h7ff1fe3;
        exp_im_rom[695] = 'h537a;
        exp_im_rom[696] = 'h7ff76fd;
        exp_im_rom[697] = 'h7ff44d1;
        exp_im_rom[698] = 'h7ff48c8;
        exp_im_rom[699] = 'h7fd1a5d;
        exp_im_rom[700] = 'h7fd92bc;
        exp_im_rom[701] = 'h7fc826e;
        exp_im_rom[702] = 'h7f84824;
        exp_im_rom[703] = 'h153984;
        exp_im_rom[704] = 'h3f497;
        exp_im_rom[705] = 'h1de35;
        exp_im_rom[706] = 'ha0a5;
        exp_im_rom[707] = 'h3a29c;
        exp_im_rom[708] = 'h135f6;
        exp_im_rom[709] = 'hae8b;
        exp_im_rom[710] = 'he3;
        exp_im_rom[711] = 'h37c5f;
        exp_im_rom[712] = 'h108b4;
        exp_im_rom[713] = 'ha170;
        exp_im_rom[714] = 'h1fe4;
        exp_im_rom[715] = 'h33c46;
        exp_im_rom[716] = 'h1198d;
        exp_im_rom[717] = 'he53a;
        exp_im_rom[718] = 'hea71;
        exp_im_rom[719] = 'h7ffaec5;
        exp_im_rom[720] = 'h7297;
        exp_im_rom[721] = 'h82c5;
        exp_im_rom[722] = 'h95c8;
        exp_im_rom[723] = 'h7fffdc5;
        exp_im_rom[724] = 'h72af;
        exp_im_rom[725] = 'h8aef;
        exp_im_rom[726] = 'hbb6a;
        exp_im_rom[727] = 'h7ff102c;
        exp_im_rom[728] = 'h6110;
        exp_im_rom[729] = 'h9911;
        exp_im_rom[730] = 'hf170;
        exp_im_rom[731] = 'h7fe54e6;
        exp_im_rom[732] = 'haff2;
        exp_im_rom[733] = 'h1696f;
        exp_im_rom[734] = 'h36a13;
        exp_im_rom[735] = 'h7e70acd;
        exp_im_rom[736] = 'h7fcef3b;
        exp_im_rom[737] = 'h7fe4ac9;
        exp_im_rom[738] = 'h7feea13;
        exp_im_rom[739] = 'h7fc0be2;
        exp_im_rom[740] = 'h7fe8b7a;
        exp_im_rom[741] = 'h7fea266;
        exp_im_rom[742] = 'h7fe660b;
        exp_im_rom[743] = 'h3d22a;
        exp_im_rom[744] = 'h7ff3e0f;
        exp_im_rom[745] = 'h7fec9fd;
        exp_im_rom[746] = 'h7fdf902;
        exp_im_rom[747] = 'hd253d;
        exp_im_rom[748] = 'h7ffcd16;
        exp_im_rom[749] = 'h7fe9dde;
        exp_im_rom[750] = 'h7fc3cde;
        exp_im_rom[751] = 'h3e2048;
        exp_im_rom[752] = 'h49a59;
        exp_im_rom[753] = 'h30953;
        exp_im_rom[754] = 'h35638;
        exp_im_rom[755] = 'h7df4f3f;
        exp_im_rom[756] = 'h7ff75b8;
        exp_im_rom[757] = 'h4ebf;
        exp_im_rom[758] = 'h110b0;
        exp_im_rom[759] = 'h7e06309;
        exp_im_rom[760] = 'h7fee989;
        exp_im_rom[761] = 'h7ff727b;
        exp_im_rom[762] = 'h7ffa36f;
        exp_im_rom[763] = 'h7fd9408;
        exp_im_rom[764] = 'h7ffa835;
        exp_im_rom[765] = 'h7ffaaca;
        exp_im_rom[766] = 'h7ff9523;
        exp_im_rom[767] = 'h343f32;
        exp_im_rom[768] = 'h7fffff8;
        exp_im_rom[769] = 'h7ffe23e;
        exp_im_rom[770] = 'h7ffce5f;
        exp_im_rom[771] = 'h7f950b9;
        exp_im_rom[772] = 'h7ffe5ee;
        exp_im_rom[773] = 'h7ffcf65;
        exp_im_rom[774] = 'h7ffad87;
        exp_im_rom[775] = 'h7f7f473;
        exp_im_rom[776] = 'he7e;
        exp_im_rom[777] = 'h7ffe4ec;
        exp_im_rom[778] = 'h7ffbbd7;
        exp_im_rom[779] = 'h7fa62ab;
        exp_im_rom[780] = 'h2756;
        exp_im_rom[781] = 'h7fffe66;
        exp_im_rom[782] = 'h7ffe4ca;
        exp_im_rom[783] = 'h7fe78c8;
        exp_im_rom[784] = 'h7fffbcf;
        exp_im_rom[785] = 'h7ffe239;
        exp_im_rom[786] = 'h7ffc23c;
        exp_im_rom[787] = 'h7fd4add;
        exp_im_rom[788] = 'h147f;
        exp_im_rom[789] = 'h7ffeaba;
        exp_im_rom[790] = 'h7ffc46d;
        exp_im_rom[791] = 'h7fda87b;
        exp_im_rom[792] = 'h1063;
        exp_im_rom[793] = 'h7ffdae9;
        exp_im_rom[794] = 'h7ff9bcd;
        exp_im_rom[795] = 'h7fc2fcd;
        exp_im_rom[796] = 'h329d;
        exp_im_rom[797] = 'h7ffb9b6;
        exp_im_rom[798] = 'h7feedfe;
        exp_im_rom[799] = 'h7f13aeb;
        exp_im_rom[800] = 'h2f2c1;
        exp_im_rom[801] = 'h21c51;
        exp_im_rom[802] = 'h297cb;
        exp_im_rom[803] = 'hf0948;
        exp_im_rom[804] = 'h7fe73a9;
        exp_im_rom[805] = 'h7ffc54d;
        exp_im_rom[806] = 'h8b9b;
        exp_im_rom[807] = 'h6ffe6;
        exp_im_rom[808] = 'h7fe890b;
        exp_im_rom[809] = 'h7ff5a6c;
        exp_im_rom[810] = 'h7ffc21a;
        exp_im_rom[811] = 'h1cc97;
        exp_im_rom[812] = 'h7ff4ada;
        exp_im_rom[813] = 'h7ffbd2d;
        exp_im_rom[814] = 'h4da2;
        exp_im_rom[815] = 'h625b0;
        exp_im_rom[816] = 'h7fdb22d;
        exp_im_rom[817] = 'h7fe8c4f;
        exp_im_rom[818] = 'h7fed726;
        exp_im_rom[819] = 'h5840;
        exp_im_rom[820] = 'h7fdd829;
        exp_im_rom[821] = 'h7fda3f8;
        exp_im_rom[822] = 'h7fc6194;
        exp_im_rom[823] = 'h7ee20fd;
        exp_im_rom[824] = 'h48f4c;
        exp_im_rom[825] = 'h22b7a;
        exp_im_rom[826] = 'h24e84;
        exp_im_rom[827] = 'hbcdfb;
        exp_im_rom[828] = 'h7fb099c;
        exp_im_rom[829] = 'h7fc4680;
        exp_im_rom[830] = 'h7fadcd1;
        exp_im_rom[831] = 'h7ea1d84;
        exp_im_rom[832] = 'h60367;
        exp_im_rom[833] = 'h1d77c;
        exp_im_rom[834] = 'h145;
        exp_im_rom[835] = 'h7f86bd1;
        exp_im_rom[836] = 'h47209;
        exp_im_rom[837] = 'h284a7;
        exp_im_rom[838] = 'h22473;
        exp_im_rom[839] = 'h3caeb;
        exp_im_rom[840] = 'h1909;
        exp_im_rom[841] = 'h82c7;
        exp_im_rom[842] = 'h84c4;
        exp_im_rom[843] = 'h2c0c;
        exp_im_rom[844] = 'hc5f8;
        exp_im_rom[845] = 'ha22f;
        exp_im_rom[846] = 'h8ae6;
        exp_im_rom[847] = 'h193f;
        exp_im_rom[848] = 'hef1b;
        exp_im_rom[849] = 'hd287;
        exp_im_rom[850] = 'he820;
        exp_im_rom[851] = 'h1d833;
        exp_im_rom[852] = 'h7ffe8e8;
        exp_im_rom[853] = 'h395c;
        exp_im_rom[854] = 'h270a;
        exp_im_rom[855] = 'h7fed2bb;
        exp_im_rom[856] = 'h1df4a;
        exp_im_rom[857] = 'h170b9;
        exp_im_rom[858] = 'h197e0;
        exp_im_rom[859] = 'h2cf40;
        exp_im_rom[860] = 'hce35;
        exp_im_rom[861] = 'h1deb4;
        exp_im_rom[862] = 'h36f2e;
        exp_im_rom[863] = 'hcc522;
        exp_im_rom[864] = 'h7f881f3;
        exp_im_rom[865] = 'h7fd3c5b;
        exp_im_rom[866] = 'h7fe929a;
        exp_im_rom[867] = 'hc432;
        exp_im_rom[868] = 'h7fcc413;
        exp_im_rom[869] = 'h7fd8fcc;
        exp_im_rom[870] = 'h7fcf197;
        exp_im_rom[871] = 'h7f6ecb7;
        exp_im_rom[872] = 'h629e5;
        exp_im_rom[873] = 'h2c56d;
        exp_im_rom[874] = 'h28d9c;
        exp_im_rom[875] = 'h4b5c6;
        exp_im_rom[876] = 'h7ffc5a8;
        exp_im_rom[877] = 'h22350;
        exp_im_rom[878] = 'h51812;
        exp_im_rom[879] = 'h151e1a;
        exp_im_rom[880] = 'h7ebc1cd;
        exp_im_rom[881] = 'h7f6c15c;
        exp_im_rom[882] = 'h7f8833b;
        exp_im_rom[883] = 'h7f727fc;
        exp_im_rom[884] = 'h7fb92f3;
        exp_im_rom[885] = 'h7f8a716;
        exp_im_rom[886] = 'h7f3fbc3;
        exp_im_rom[887] = 'h7dadecd;
        exp_im_rom[888] = 'h2153b8;
        exp_im_rom[889] = 'hcea2e;
        exp_im_rom[890] = 'ha8502;
        exp_im_rom[891] = 'h13c62d;
        exp_im_rom[892] = 'h7f1735b;
        exp_im_rom[893] = 'h7fa4931;
        exp_im_rom[894] = 'h7f9badb;
        exp_im_rom[895] = 'h7eeb5e6;
        exp_im_rom[896] = 'h122679;
        exp_im_rom[897] = 'h6ea1a;
        exp_im_rom[898] = 'h51c0f;
        exp_im_rom[899] = 'h5e2a2;
        exp_im_rom[900] = 'hd845;
        exp_im_rom[901] = 'h2aef0;
        exp_im_rom[902] = 'h3f591;
        exp_im_rom[903] = 'h99526;
        exp_im_rom[904] = 'h7f72228;
        exp_im_rom[905] = 'h7fdb04f;
        exp_im_rom[906] = 'h7fee06e;
        exp_im_rom[907] = 'h7ff43ac;
        exp_im_rom[908] = 'h7ffd9da;
        exp_im_rom[909] = 'h7ffde52;
        exp_im_rom[910] = 'h7ffed1c;
        exp_im_rom[911] = 'h7ffec33;
        exp_im_rom[912] = 'h1e8e;
        exp_im_rom[913] = 'hc5e;
        exp_im_rom[914] = 'h7fffcbb;
        exp_im_rom[915] = 'h7ffbef0;
        exp_im_rom[916] = 'h6f83;
        exp_im_rom[917] = 'h7ffefa0;
        exp_im_rom[918] = 'h7ff5d9e;
        exp_im_rom[919] = 'h7fcbcac;
        exp_im_rom[920] = 'h7b2ac;
        exp_im_rom[921] = 'h3816f;
        exp_im_rom[922] = 'h36aaf;
        exp_im_rom[923] = 'h5ab92;
        exp_im_rom[924] = 'h7fbf065;
        exp_im_rom[925] = 'h9b27;
        exp_im_rom[926] = 'h2555b;
        exp_im_rom[927] = 'h743f0;
        exp_im_rom[928] = 'h7f2dd4e;
        exp_im_rom[929] = 'h7fc10a9;
        exp_im_rom[930] = 'h7fd483a;
        exp_im_rom[931] = 'h7fcb07b;
        exp_im_rom[932] = 'h28ac8;
        exp_im_rom[933] = 'h1e04;
        exp_im_rom[934] = 'h7ffb637;
        exp_im_rom[935] = 'h7fece4e;
        exp_im_rom[936] = 'h39702;
        exp_im_rom[937] = 'h19e88;
        exp_im_rom[938] = 'h1dc63;
        exp_im_rom[939] = 'h3ceb0;
        exp_im_rom[940] = 'h7f9e861;
        exp_im_rom[941] = 'h7ff3048;
        exp_im_rom[942] = 'h810f;
        exp_im_rom[943] = 'h3508a;
        exp_im_rom[944] = 'h7f56752;
        exp_im_rom[945] = 'h7fca1ca;
        exp_im_rom[946] = 'h7fd5a08;
        exp_im_rom[947] = 'h7fc914f;
        exp_im_rom[948] = 'h387fd;
        exp_im_rom[949] = 'h7ffec2f;
        exp_im_rom[950] = 'h7ff56d9;
        exp_im_rom[951] = 'h7fe7454;
        exp_im_rom[952] = 'h2be7e;
        exp_im_rom[953] = 'h4cb;
        exp_im_rom[954] = 'h7ff1599;
        exp_im_rom[955] = 'h7fc28c9;
        exp_im_rom[956] = 'h10b417;
        exp_im_rom[957] = 'h5c759;
        exp_im_rom[958] = 'h60d48;
        exp_im_rom[959] = 'hba3a4;
        exp_im_rom[960] = 'h7e08474;
        exp_im_rom[961] = 'h7f9ef43;
        exp_im_rom[962] = 'h7fc9545;
        exp_im_rom[963] = 'h7fd3cb6;
        exp_im_rom[964] = 'hb6a6;
        exp_im_rom[965] = 'h7ff4f88;
        exp_im_rom[966] = 'h7ff866e;
        exp_im_rom[967] = 'h5605;
        exp_im_rom[968] = 'h7fa4a13;
        exp_im_rom[969] = 'h7fe3a50;
        exp_im_rom[970] = 'h7fea00d;
        exp_im_rom[971] = 'h7feb4eb;
        exp_im_rom[972] = 'h7ffa17f;
        exp_im_rom[973] = 'h7ff25a4;
        exp_im_rom[974] = 'h7ff23cc;
        exp_im_rom[975] = 'h7ff2906;
        exp_im_rom[976] = 'h7fefb17;
        exp_im_rom[977] = 'h7ff15fd;
        exp_im_rom[978] = 'h7ff0e8e;
        exp_im_rom[979] = 'h7fef0ab;
        exp_im_rom[980] = 'h7fff1e8;
        exp_im_rom[981] = 'h7ff2458;
        exp_im_rom[982] = 'h7fef1e1;
        exp_im_rom[983] = 'h7fe7d7a;
        exp_im_rom[984] = 'h32f5c;
        exp_im_rom[985] = 'h7ffa5b7;
        exp_im_rom[986] = 'h7ff44f2;
        exp_im_rom[987] = 'h7fedaf3;
        exp_im_rom[988] = 'h1fd49;
        exp_im_rom[989] = 'h7ff4e65;
        exp_im_rom[990] = 'h7fec3aa;
        exp_im_rom[991] = 'h7fd8bd1;
        exp_im_rom[992] = 'he2035;
        exp_im_rom[993] = 'h11517;
        exp_im_rom[994] = 'h29f0;
        exp_im_rom[995] = 'h7ff78b6;
        exp_im_rom[996] = 'h5c6a4;
        exp_im_rom[997] = 'h6802;
        exp_im_rom[998] = 'h7fff1ec;
        exp_im_rom[999] = 'h7ff6d39;
        exp_im_rom[1000] = 'h67b25;
        exp_im_rom[1001] = 'h6fd5;
        exp_im_rom[1002] = 'h84f;
        exp_im_rom[1003] = 'h7ffa0da;
        exp_im_rom[1004] = 'h5dc11;
        exp_im_rom[1005] = 'h595a;
        exp_im_rom[1006] = 'h34a;
        exp_im_rom[1007] = 'h7ff9f61;
        exp_im_rom[1008] = 'h85290;
        exp_im_rom[1009] = 'h8910;
        exp_im_rom[1010] = 'h3e1d;
        exp_im_rom[1011] = 'hed4;
        exp_im_rom[1012] = 'h31c22;
        exp_im_rom[1013] = 'h38ce;
        exp_im_rom[1014] = 'h1bbe;
        exp_im_rom[1015] = 'h26b;
        exp_im_rom[1016] = 'h33794;
        exp_im_rom[1017] = 'h267f;
        exp_im_rom[1018] = 'h1503;
        exp_im_rom[1019] = 'ha54;
        exp_im_rom[1020] = 'h149b0;
        exp_im_rom[1021] = 'hb28;
        exp_im_rom[1022] = 'h5c7;
        exp_im_rom[1023] = 'h284;
    end
    else begin
        exp_im_rom[0] = 'h7fffeaa;
        exp_im_rom[1] = 'h243;
        exp_im_rom[2] = 'h5aa;
        exp_im_rom[3] = 'hb31;
        exp_im_rom[4] = 'h149b0;
        exp_im_rom[5] = 'ha67;
        exp_im_rom[6] = 'h14e2;
        exp_im_rom[7] = 'h266e;
        exp_im_rom[8] = 'h33793;
        exp_im_rom[9] = 'h27c;
        exp_im_rom[10] = 'h1bc8;
        exp_im_rom[11] = 'h38d6;
        exp_im_rom[12] = 'h31c26;
        exp_im_rom[13] = 'hee4;
        exp_im_rom[14] = 'h3e1f;
        exp_im_rom[15] = 'h890b;
        exp_im_rom[16] = 'h85296;
        exp_im_rom[17] = 'h7ff9f95;
        exp_im_rom[18] = 'h356;
        exp_im_rom[19] = 'h5954;
        exp_im_rom[20] = 'h5dc0d;
        exp_im_rom[21] = 'h7ffa0cd;
        exp_im_rom[22] = 'h85a;
        exp_im_rom[23] = 'h6fdb;
        exp_im_rom[24] = 'h67b2e;
        exp_im_rom[25] = 'h7ff6d55;
        exp_im_rom[26] = 'h7fff1e6;
        exp_im_rom[27] = 'h67fd;
        exp_im_rom[28] = 'h5c69a;
        exp_im_rom[29] = 'h7ff78a7;
        exp_im_rom[30] = 'h2a09;
        exp_im_rom[31] = 'h114e0;
        exp_im_rom[32] = 'he202e;
        exp_im_rom[33] = 'h7fd8be5;
        exp_im_rom[34] = 'h7fec38a;
        exp_im_rom[35] = 'h7ff4e55;
        exp_im_rom[36] = 'h1fd49;
        exp_im_rom[37] = 'h7fedaf7;
        exp_im_rom[38] = 'h7ff44d4;
        exp_im_rom[39] = 'h7ffa5ab;
        exp_im_rom[40] = 'h32f68;
        exp_im_rom[41] = 'h7fe7d56;
        exp_im_rom[42] = 'h7fef1d7;
        exp_im_rom[43] = 'h7ff2453;
        exp_im_rom[44] = 'h7fff1ed;
        exp_im_rom[45] = 'h7fef0a4;
        exp_im_rom[46] = 'h7ff0e92;
        exp_im_rom[47] = 'h7ff1604;
        exp_im_rom[48] = 'h7fefb16;
        exp_im_rom[49] = 'h7ff2900;
        exp_im_rom[50] = 'h7ff23bf;
        exp_im_rom[51] = 'h7ff25af;
        exp_im_rom[52] = 'h7ffa178;
        exp_im_rom[53] = 'h7feb4e3;
        exp_im_rom[54] = 'h7fea012;
        exp_im_rom[55] = 'h7fe3a5e;
        exp_im_rom[56] = 'h7fa4a0b;
        exp_im_rom[57] = 'h5615;
        exp_im_rom[58] = 'h7ff8663;
        exp_im_rom[59] = 'h7ff4f85;
        exp_im_rom[60] = 'hb6a3;
        exp_im_rom[61] = 'h7fd3cbc;
        exp_im_rom[62] = 'h7fc9547;
        exp_im_rom[63] = 'h7f9ef2a;
        exp_im_rom[64] = 'h7e08474;
        exp_im_rom[65] = 'hba3d3;
        exp_im_rom[66] = 'h60d74;
        exp_im_rom[67] = 'h5c754;
        exp_im_rom[68] = 'h10b424;
        exp_im_rom[69] = 'h7fc28d4;
        exp_im_rom[70] = 'h7ff1590;
        exp_im_rom[71] = 'h4c9;
        exp_im_rom[72] = 'h2be7c;
        exp_im_rom[73] = 'h7fe7456;
        exp_im_rom[74] = 'h7ff56ea;
        exp_im_rom[75] = 'h7ffec33;
        exp_im_rom[76] = 'h38803;
        exp_im_rom[77] = 'h7fc9152;
        exp_im_rom[78] = 'h7fd5a23;
        exp_im_rom[79] = 'h7fca1ad;
        exp_im_rom[80] = 'h7f56747;
        exp_im_rom[81] = 'h35088;
        exp_im_rom[82] = 'h80fc;
        exp_im_rom[83] = 'h7ff304b;
        exp_im_rom[84] = 'h7f9e854;
        exp_im_rom[85] = 'h3ceb4;
        exp_im_rom[86] = 'h1dc6f;
        exp_im_rom[87] = 'h19e98;
        exp_im_rom[88] = 'h396f9;
        exp_im_rom[89] = 'h7fece4b;
        exp_im_rom[90] = 'h7ffb649;
        exp_im_rom[91] = 'h1e09;
        exp_im_rom[92] = 'h28abf;
        exp_im_rom[93] = 'h7fcb08d;
        exp_im_rom[94] = 'h7fd4820;
        exp_im_rom[95] = 'h7fc109e;
        exp_im_rom[96] = 'h7f2dd42;
        exp_im_rom[97] = 'h743e4;
        exp_im_rom[98] = 'h2553a;
        exp_im_rom[99] = 'h9b39;
        exp_im_rom[100] = 'h7fbf061;
        exp_im_rom[101] = 'h5ab8e;
        exp_im_rom[102] = 'h36aa4;
        exp_im_rom[103] = 'h3818f;
        exp_im_rom[104] = 'h7b2b5;
        exp_im_rom[105] = 'h7fcbca6;
        exp_im_rom[106] = 'h7ff5da2;
        exp_im_rom[107] = 'h7ffef9f;
        exp_im_rom[108] = 'h6f81;
        exp_im_rom[109] = 'h7ffbef3;
        exp_im_rom[110] = 'h7fffcdc;
        exp_im_rom[111] = 'hc51;
        exp_im_rom[112] = 'h1e94;
        exp_im_rom[113] = 'h7ffec61;
        exp_im_rom[114] = 'h7ffed1d;
        exp_im_rom[115] = 'h7ffde5b;
        exp_im_rom[116] = 'h7ffd9d9;
        exp_im_rom[117] = 'h7ff439d;
        exp_im_rom[118] = 'h7fee076;
        exp_im_rom[119] = 'h7fdb065;
        exp_im_rom[120] = 'h7f72228;
        exp_im_rom[121] = 'h9952b;
        exp_im_rom[122] = 'h3f5a3;
        exp_im_rom[123] = 'h2aef6;
        exp_im_rom[124] = 'hd84f;
        exp_im_rom[125] = 'h5e2ad;
        exp_im_rom[126] = 'h51c1b;
        exp_im_rom[127] = 'h6ea2a;
        exp_im_rom[128] = 'h122679;
        exp_im_rom[129] = 'h7eeb61e;
        exp_im_rom[130] = 'h7f9bacd;
        exp_im_rom[131] = 'h7fa492e;
        exp_im_rom[132] = 'h7f17358;
        exp_im_rom[133] = 'h13c614;
        exp_im_rom[134] = 'ha84d7;
        exp_im_rom[135] = 'hcea28;
        exp_im_rom[136] = 'h2153ac;
        exp_im_rom[137] = 'h7dadee5;
        exp_im_rom[138] = 'h7f3fbe5;
        exp_im_rom[139] = 'h7f8a717;
        exp_im_rom[140] = 'h7fb92f7;
        exp_im_rom[141] = 'h7f727e3;
        exp_im_rom[142] = 'h7f88366;
        exp_im_rom[143] = 'h7f6c15c;
        exp_im_rom[144] = 'h7ebc1e3;
        exp_im_rom[145] = 'h151dfd;
        exp_im_rom[146] = 'h517ed;
        exp_im_rom[147] = 'h2234a;
        exp_im_rom[148] = 'h7ffc5ad;
        exp_im_rom[149] = 'h4b5d1;
        exp_im_rom[150] = 'h28d83;
        exp_im_rom[151] = 'h2c57a;
        exp_im_rom[152] = 'h629df;
        exp_im_rom[153] = 'h7f6ecb0;
        exp_im_rom[154] = 'h7fcf175;
        exp_im_rom[155] = 'h7fd8fde;
        exp_im_rom[156] = 'h7fcc422;
        exp_im_rom[157] = 'hc42e;
        exp_im_rom[158] = 'h7fe928d;
        exp_im_rom[159] = 'h7fd3c8c;
        exp_im_rom[160] = 'h7f88209;
        exp_im_rom[161] = 'hcc50d;
        exp_im_rom[162] = 'h36f13;
        exp_im_rom[163] = 'h1debe;
        exp_im_rom[164] = 'hce33;
        exp_im_rom[165] = 'h2cf38;
        exp_im_rom[166] = 'h197df;
        exp_im_rom[167] = 'h170ae;
        exp_im_rom[168] = 'h1df50;
        exp_im_rom[169] = 'h7fed2c5;
        exp_im_rom[170] = 'h2724;
        exp_im_rom[171] = 'h3951;
        exp_im_rom[172] = 'h7ffe8e3;
        exp_im_rom[173] = 'h1d830;
        exp_im_rom[174] = 'he847;
        exp_im_rom[175] = 'hd285;
        exp_im_rom[176] = 'hef1b;
        exp_im_rom[177] = 'h193f;
        exp_im_rom[178] = 'h8aee;
        exp_im_rom[179] = 'ha224;
        exp_im_rom[180] = 'hc5f0;
        exp_im_rom[181] = 'h2c02;
        exp_im_rom[182] = 'h84d7;
        exp_im_rom[183] = 'h82ce;
        exp_im_rom[184] = 'h18fd;
        exp_im_rom[185] = 'h3caeb;
        exp_im_rom[186] = 'h2246d;
        exp_im_rom[187] = 'h284b6;
        exp_im_rom[188] = 'h47217;
        exp_im_rom[189] = 'h7f86be2;
        exp_im_rom[190] = 'h12c;
        exp_im_rom[191] = 'h1d795;
        exp_im_rom[192] = 'h60367;
        exp_im_rom[193] = 'h7ea1d61;
        exp_im_rom[194] = 'h7fadcdd;
        exp_im_rom[195] = 'h7fc46a0;
        exp_im_rom[196] = 'h7fb09a9;
        exp_im_rom[197] = 'hbce08;
        exp_im_rom[198] = 'h24e7f;
        exp_im_rom[199] = 'h22b6a;
        exp_im_rom[200] = 'h48f3e;
        exp_im_rom[201] = 'h7ee2105;
        exp_im_rom[202] = 'h7fc618e;
        exp_im_rom[203] = 'h7fda3ff;
        exp_im_rom[204] = 'h7fdd831;
        exp_im_rom[205] = 'h5843;
        exp_im_rom[206] = 'h7fed738;
        exp_im_rom[207] = 'h7fe8c54;
        exp_im_rom[208] = 'h7fdb22f;
        exp_im_rom[209] = 'h625a4;
        exp_im_rom[210] = 'h4da9;
        exp_im_rom[211] = 'h7ffbd19;
        exp_im_rom[212] = 'h7ff4adc;
        exp_im_rom[213] = 'h1cc98;
        exp_im_rom[214] = 'h7ffc214;
        exp_im_rom[215] = 'h7ff5a6f;
        exp_im_rom[216] = 'h7fe8903;
        exp_im_rom[217] = 'h6ffe0;
        exp_im_rom[218] = 'h8ba5;
        exp_im_rom[219] = 'h7ffc551;
        exp_im_rom[220] = 'h7fe73ad;
        exp_im_rom[221] = 'hf0958;
        exp_im_rom[222] = 'h297f9;
        exp_im_rom[223] = 'h21c65;
        exp_im_rom[224] = 'h2f2c5;
        exp_im_rom[225] = 'h7f13aed;
        exp_im_rom[226] = 'h7feee06;
        exp_im_rom[227] = 'h7ffb9b1;
        exp_im_rom[228] = 'h32a4;
        exp_im_rom[229] = 'h7fc2fbb;
        exp_im_rom[230] = 'h7ff9bd4;
        exp_im_rom[231] = 'h7ffdade;
        exp_im_rom[232] = 'h105b;
        exp_im_rom[233] = 'h7fda865;
        exp_im_rom[234] = 'h7ffc455;
        exp_im_rom[235] = 'h7ffeaba;
        exp_im_rom[236] = 'h1485;
        exp_im_rom[237] = 'h7fd4ad5;
        exp_im_rom[238] = 'h7ffc23f;
        exp_im_rom[239] = 'h7ffe249;
        exp_im_rom[240] = 'h7fffbd2;
        exp_im_rom[241] = 'h7fe78d0;
        exp_im_rom[242] = 'h7ffe4de;
        exp_im_rom[243] = 'h7fffe50;
        exp_im_rom[244] = 'h2759;
        exp_im_rom[245] = 'h7fa62b3;
        exp_im_rom[246] = 'h7ffbbc8;
        exp_im_rom[247] = 'h7ffe4fa;
        exp_im_rom[248] = 'he79;
        exp_im_rom[249] = 'h7f7f46f;
        exp_im_rom[250] = 'h7ffadaf;
        exp_im_rom[251] = 'h7ffcf70;
        exp_im_rom[252] = 'h7ffe5e8;
        exp_im_rom[253] = 'h7f950bd;
        exp_im_rom[254] = 'h7ffce61;
        exp_im_rom[255] = 'h7ffe25a;
        exp_im_rom[256] = 'h7fffff8;
        exp_im_rom[257] = 'h343f19;
        exp_im_rom[258] = 'h7ff954a;
        exp_im_rom[259] = 'h7ffaada;
        exp_im_rom[260] = 'h7ffa837;
        exp_im_rom[261] = 'h7fd93fa;
        exp_im_rom[262] = 'h7ffa37d;
        exp_im_rom[263] = 'h7ff728f;
        exp_im_rom[264] = 'h7fee98d;
        exp_im_rom[265] = 'h7e0630c;
        exp_im_rom[266] = 'h110be;
        exp_im_rom[267] = 'h4ebd;
        exp_im_rom[268] = 'h7ff75b8;
        exp_im_rom[269] = 'h7df4f37;
        exp_im_rom[270] = 'h3562e;
        exp_im_rom[271] = 'h30938;
        exp_im_rom[272] = 'h49a52;
        exp_im_rom[273] = 'h3e2042;
        exp_im_rom[274] = 'h7fc3cf7;
        exp_im_rom[275] = 'h7fe9dd2;
        exp_im_rom[276] = 'h7ffcd0e;
        exp_im_rom[277] = 'hd2550;
        exp_im_rom[278] = 'h7fdf8f4;
        exp_im_rom[279] = 'h7fec9f1;
        exp_im_rom[280] = 'h7ff3e16;
        exp_im_rom[281] = 'h3d226;
        exp_im_rom[282] = 'h7fe6616;
        exp_im_rom[283] = 'h7fea267;
        exp_im_rom[284] = 'h7fe8b80;
        exp_im_rom[285] = 'h7fc0bc4;
        exp_im_rom[286] = 'h7feea2a;
        exp_im_rom[287] = 'h7fe4aba;
        exp_im_rom[288] = 'h7fcef37;
        exp_im_rom[289] = 'h7e70ada;
        exp_im_rom[290] = 'h36a28;
        exp_im_rom[291] = 'h16976;
        exp_im_rom[292] = 'hafe4;
        exp_im_rom[293] = 'h7fe54d7;
        exp_im_rom[294] = 'hf169;
        exp_im_rom[295] = 'h9911;
        exp_im_rom[296] = 'h6101;
        exp_im_rom[297] = 'h7ff1026;
        exp_im_rom[298] = 'hbb6a;
        exp_im_rom[299] = 'h8ae3;
        exp_im_rom[300] = 'h72ab;
        exp_im_rom[301] = 'h7fffdc6;
        exp_im_rom[302] = 'h95d8;
        exp_im_rom[303] = 'h82c5;
        exp_im_rom[304] = 'h7296;
        exp_im_rom[305] = 'h7ffaee0;
        exp_im_rom[306] = 'hea6e;
        exp_im_rom[307] = 'he532;
        exp_im_rom[308] = 'h11996;
        exp_im_rom[309] = 'h33c3e;
        exp_im_rom[310] = 'h1fd6;
        exp_im_rom[311] = 'ha160;
        exp_im_rom[312] = 'h108b8;
        exp_im_rom[313] = 'h37c5b;
        exp_im_rom[314] = 'h101;
        exp_im_rom[315] = 'hae93;
        exp_im_rom[316] = 'h13605;
        exp_im_rom[317] = 'h3a2bc;
        exp_im_rom[318] = 'ha098;
        exp_im_rom[319] = 'h1de36;
        exp_im_rom[320] = 'h3f497;
        exp_im_rom[321] = 'h153989;
        exp_im_rom[322] = 'h7f847f3;
        exp_im_rom[323] = 'h7fc8248;
        exp_im_rom[324] = 'h7fd92c6;
        exp_im_rom[325] = 'h7fd1a70;
        exp_im_rom[326] = 'h7ff48bc;
        exp_im_rom[327] = 'h7ff44ca;
        exp_im_rom[328] = 'h7ff7712;
        exp_im_rom[329] = 'h5382;
        exp_im_rom[330] = 'h7ff1fde;
        exp_im_rom[331] = 'h7ff876a;
        exp_im_rom[332] = 'h7fff193;
        exp_im_rom[333] = 'h249ad;
        exp_im_rom[334] = 'h7fe2a5a;
        exp_im_rom[335] = 'h7ff0797;
        exp_im_rom[336] = 'h7ff77f9;
        exp_im_rom[337] = 'h14777;
        exp_im_rom[338] = 'h7fdf4fc;
        exp_im_rom[339] = 'h7fe8945;
        exp_im_rom[340] = 'h7fe7a61;
        exp_im_rom[341] = 'h7fcc6c2;
        exp_im_rom[342] = 'h73a5;
        exp_im_rom[343] = 'h7ffc67d;
        exp_im_rom[344] = 'h7ffa149;
        exp_im_rom[345] = 'h7ffa023;
        exp_im_rom[346] = 'h7ff6c49;
        exp_im_rom[347] = 'h7ff5d1f;
        exp_im_rom[348] = 'h7ff25b1;
        exp_im_rom[349] = 'h7fd92ae;
        exp_im_rom[350] = 'h11f76;
        exp_im_rom[351] = 'h7a8d;
        exp_im_rom[352] = 'h9e21;
        exp_im_rom[353] = 'h29fd5;
        exp_im_rom[354] = 'h7fdd720;
        exp_im_rom[355] = 'h7fed7d9;
        exp_im_rom[356] = 'h7fee6dd;
        exp_im_rom[357] = 'h7fde270;
        exp_im_rom[358] = 'h8751;
        exp_im_rom[359] = 'h7ffe943;
        exp_im_rom[360] = 'h7ffbeb5;
        exp_im_rom[361] = 'h7ff683b;
        exp_im_rom[362] = 'h1bff;
        exp_im_rom[363] = 'h7ffeae9;
        exp_im_rom[364] = 'h7ffdd93;
        exp_im_rom[365] = 'h7ffbe21;
        exp_im_rom[366] = 'h116f;
        exp_im_rom[367] = 'h540;
        exp_im_rom[368] = 'h1394;
        exp_im_rom[369] = 'h66bd;
        exp_im_rom[370] = 'h7ff9f22;
        exp_im_rom[371] = 'h7ffde52;
        exp_im_rom[372] = 'h7ffe48a;
        exp_im_rom[373] = 'h7ff6287;
        exp_im_rom[374] = 'h17140;
        exp_im_rom[375] = 'h14d33;
        exp_im_rom[376] = 'h210a0;
        exp_im_rom[377] = 'h63a6b;
        exp_im_rom[378] = 'h7fb1649;
        exp_im_rom[379] = 'h7ff24c6;
        exp_im_rom[380] = 'h13f8a;
        exp_im_rom[381] = 'h93ddb;
        exp_im_rom[382] = 'h7f1b899;
        exp_im_rom[383] = 'h7f893b6;
        exp_im_rom[384] = 'h7f842b1;
        exp_im_rom[385] = 'h7ef225e;
        exp_im_rom[386] = 'he2b47;
        exp_im_rom[387] = 'h48f41;
        exp_im_rom[388] = 'h3b71f;
        exp_im_rom[389] = 'h80116;
        exp_im_rom[390] = 'h7f76a63;
        exp_im_rom[391] = 'h7fcc638;
        exp_im_rom[392] = 'h7fd8095;
        exp_im_rom[393] = 'h7fce405;
        exp_im_rom[394] = 'h3e87;
        exp_im_rom[395] = 'h7ff347c;
        exp_im_rom[396] = 'h7ff3270;
        exp_im_rom[397] = 'h3994;
        exp_im_rom[398] = 'h7fb9544;
        exp_im_rom[399] = 'h7fcc510;
        exp_im_rom[400] = 'h7fc0651;
        exp_im_rom[401] = 'h7f774aa;
        exp_im_rom[402] = 'h8be24;
        exp_im_rom[403] = 'h2324e;
        exp_im_rom[404] = 'h1c0d5;
        exp_im_rom[405] = 'h59d60;
        exp_im_rom[406] = 'h7f1e7ee;
        exp_im_rom[407] = 'h7f7e875;
        exp_im_rom[408] = 'h7f5af84;
        exp_im_rom[409] = 'h7e7380b;
        exp_im_rom[410] = 'h233095;
        exp_im_rom[411] = 'h9a1d2;
        exp_im_rom[412] = 'h52050;
        exp_im_rom[413] = 'h1809b;
        exp_im_rom[414] = 'ha365a;
        exp_im_rom[415] = 'h63d92;
        exp_im_rom[416] = 'h6b8a4;
        exp_im_rom[417] = 'hc7620;
        exp_im_rom[418] = 'h7f07c31;
        exp_im_rom[419] = 'h7fd14a7;
        exp_im_rom[420] = 'h7ff0be7;
        exp_im_rom[421] = 'h55cb;
        exp_im_rom[422] = 'h7fdf4ec;
        exp_im_rom[423] = 'h7ff927a;
        exp_im_rom[424] = 'h2637;
        exp_im_rom[425] = 'h16a48;
        exp_im_rom[426] = 'h7fbf701;
        exp_im_rom[427] = 'h7fec5b9;
        exp_im_rom[428] = 'h7ff3c28;
        exp_im_rom[429] = 'h7ff8fc0;
        exp_im_rom[430] = 'h7fedfe9;
        exp_im_rom[431] = 'h7ff56c0;
        exp_im_rom[432] = 'h7ff7219;
        exp_im_rom[433] = 'h7ff8f27;
        exp_im_rom[434] = 'h7ff299d;
        exp_im_rom[435] = 'h7ff608c;
        exp_im_rom[436] = 'h7ff5cb4;
        exp_im_rom[437] = 'h7ff1f69;
        exp_im_rom[438] = 'hf57e;
        exp_im_rom[439] = 'h2816;
        exp_im_rom[440] = 'h70b8;
        exp_im_rom[441] = 'h22873;
        exp_im_rom[442] = 'h7f5e551;
        exp_im_rom[443] = 'h7fc5c66;
        exp_im_rom[444] = 'h7fc73ae;
        exp_im_rom[445] = 'h7fa4c1b;
        exp_im_rom[446] = 'h9f072;
        exp_im_rom[447] = 'h6cc5;
        exp_im_rom[448] = 'h7fe9be4;
        exp_im_rom[449] = 'h7fb2ba8;
        exp_im_rom[450] = 'h119eb1;
        exp_im_rom[451] = 'h3e528;
        exp_im_rom[452] = 'h2974b;
        exp_im_rom[453] = 'h2e7c4;
        exp_im_rom[454] = 'h7fb18c5;
        exp_im_rom[455] = 'h7ff7a25;
        exp_im_rom[456] = 'h7ff9575;
        exp_im_rom[457] = 'h7feaf0e;
        exp_im_rom[458] = 'h83efb;
        exp_im_rom[459] = 'h28c5f;
        exp_im_rom[460] = 'h2cc0f;
        exp_im_rom[461] = 'h5a0c2;
        exp_im_rom[462] = 'h7e88114;
        exp_im_rom[463] = 'h7fbaa24;
        exp_im_rom[464] = 'h7fcffab;
        exp_im_rom[465] = 'h7fc7a62;
        exp_im_rom[466] = 'h80152;
        exp_im_rom[467] = 'h6cec;
        exp_im_rom[468] = 'h9a1;
        exp_im_rom[469] = 'h926b;
        exp_im_rom[470] = 'h7f7170e;
        exp_im_rom[471] = 'h7fd64dd;
        exp_im_rom[472] = 'h7fd602d;
        exp_im_rom[473] = 'h7fc276b;
        exp_im_rom[474] = 'haa27a;
        exp_im_rom[475] = 'h7ff3e69;
        exp_im_rom[476] = 'h7fd62c0;
        exp_im_rom[477] = 'h7f95b04;
        exp_im_rom[478] = 'h2e52e3;
        exp_im_rom[479] = 'h5b0a6;
        exp_im_rom[480] = 'h328cc;
        exp_im_rom[481] = 'h260d2;
        exp_im_rom[482] = 'h7ff3930;
        exp_im_rom[483] = 'h1058a;
        exp_im_rom[484] = 'hef91;
        exp_im_rom[485] = 'hd54e;
        exp_im_rom[486] = 'hd8af;
        exp_im_rom[487] = 'hbb65;
        exp_im_rom[488] = 'hbcb5;
        exp_im_rom[489] = 'heaed;
        exp_im_rom[490] = 'h7fba15c;
        exp_im_rom[491] = 'h143;
        exp_im_rom[492] = 'h2b88;
        exp_im_rom[493] = 'h4710;
        exp_im_rom[494] = 'h7fdedd9;
        exp_im_rom[495] = 'h7ffee95;
        exp_im_rom[496] = 'h7fff447;
        exp_im_rom[497] = 'h7ffdf60;
        exp_im_rom[498] = 'h29beb;
        exp_im_rom[499] = 'h17ce;
        exp_im_rom[500] = 'h7fff275;
        exp_im_rom[501] = 'h7ffb4eb;
        exp_im_rom[502] = 'h9826b;
        exp_im_rom[503] = 'h5d95;
        exp_im_rom[504] = 'h1ecc;
        exp_im_rom[505] = 'h7ffe33e;
        exp_im_rom[506] = 'hc6e3b;
        exp_im_rom[507] = 'h5b6b;
        exp_im_rom[508] = 'h2685;
        exp_im_rom[509] = 'h7fff7c8;
        exp_im_rom[510] = 'h191499;
        exp_im_rom[511] = 'h372a;
        exp_im_rom[512] = 'h6;
        exp_im_rom[513] = 'h7ffaad5;
        exp_im_rom[514] = 'h7ba8732;
        exp_im_rom[515] = 'ha331;
        exp_im_rom[516] = 'h3e5e;
        exp_im_rom[517] = 'h7ffd23f;
        exp_im_rom[518] = 'h7e3a89c;
        exp_im_rom[519] = 'h118e6;
        exp_im_rom[520] = 'hb74d;
        exp_im_rom[521] = 'h880e;
        exp_im_rom[522] = 'h7fcc552;
        exp_im_rom[523] = 'hc0fc;
        exp_im_rom[524] = 'ha244;
        exp_im_rom[525] = 'h71e2;
        exp_im_rom[526] = 'h7f7838f;
        exp_im_rom[527] = 'h1d179;
        exp_im_rom[528] = 'h1f048;
        exp_im_rom[529] = 'h2f4dd;
        exp_im_rom[530] = 'h2199c8;
        exp_im_rom[531] = 'h7fe82f0;
        exp_im_rom[532] = 'h1809;
        exp_im_rom[533] = 'h149af;
        exp_im_rom[534] = 'h128632;
        exp_im_rom[535] = 'h7fed1f9;
        exp_im_rom[536] = 'h50a0;
        exp_im_rom[537] = 'h213b5;
        exp_im_rom[538] = 'h1e9b44;
        exp_im_rom[539] = 'h7fc464d;
        exp_im_rom[540] = 'h7feb68a;
        exp_im_rom[541] = 'hf5d5;
        exp_im_rom[542] = 'h21bd0b;
        exp_im_rom[543] = 'h7f7fb46;
        exp_im_rom[544] = 'h7f9d11a;
        exp_im_rom[545] = 'h7f849eb;
        exp_im_rom[546] = 'h7d29c92;
        exp_im_rom[547] = 'h49e37;
        exp_im_rom[548] = 'h11e4d;
        exp_im_rom[549] = 'h7ffd6c9;
        exp_im_rom[550] = 'h7fac862;
        exp_im_rom[551] = 'hbb75;
        exp_im_rom[552] = 'h7ffffea;
        exp_im_rom[553] = 'h7ff821c;
        exp_im_rom[554] = 'h7fc1fb5;
        exp_im_rom[555] = 'h8caf;
        exp_im_rom[556] = 'h1201;
        exp_im_rom[557] = 'h7ffe30c;
        exp_im_rom[558] = 'h7ffb140;
        exp_im_rom[559] = 'h7ffbee4;
        exp_im_rom[560] = 'h7ffab98;
        exp_im_rom[561] = 'h7ff9b7a;
        exp_im_rom[562] = 'h7ff7377;
        exp_im_rom[563] = 'h7ff9505;
        exp_im_rom[564] = 'h7ff8a96;
        exp_im_rom[565] = 'h7ff8fc9;
        exp_im_rom[566] = 'h5f28;
        exp_im_rom[567] = 'h7feeea2;
        exp_im_rom[568] = 'h7fef6a9;
        exp_im_rom[569] = 'h7febb91;
        exp_im_rom[570] = 'h7fc50b3;
        exp_im_rom[571] = 'h3327;
        exp_im_rom[572] = 'h7ffd6f9;
        exp_im_rom[573] = 'h42dc;
        exp_im_rom[574] = 'h71e15;
        exp_im_rom[575] = 'h7faaf1e;
        exp_im_rom[576] = 'h7fb66ee;
        exp_im_rom[577] = 'h7f9994d;
        exp_im_rom[578] = 'h7e70c44;
        exp_im_rom[579] = 'h686fa;
        exp_im_rom[580] = 'h18048;
        exp_im_rom[581] = 'h7ff4e1a;
        exp_im_rom[582] = 'h7f7056e;
        exp_im_rom[583] = 'h41351;
        exp_im_rom[584] = 'h196be;
        exp_im_rom[585] = 'h9656;
        exp_im_rom[586] = 'h7fe6f42;
        exp_im_rom[587] = 'h11359;
        exp_im_rom[588] = 'h178f;
        exp_im_rom[589] = 'h7ff189c;
        exp_im_rom[590] = 'h7f98fd9;
        exp_im_rom[591] = 'h36e3b;
        exp_im_rom[592] = 'h17087;
        exp_im_rom[593] = 'hb72a;
        exp_im_rom[594] = 'h7ff6148;
        exp_im_rom[595] = 'h1079b;
        exp_im_rom[596] = 'h56a6;
        exp_im_rom[597] = 'h7ffac1e;
        exp_im_rom[598] = 'h7fc57c1;
        exp_im_rom[599] = 'h2a540;
        exp_im_rom[600] = 'h135d7;
        exp_im_rom[601] = 'hb393;
        exp_im_rom[602] = 'h7ffdfa9;
        exp_im_rom[603] = 'hcda1;
        exp_im_rom[604] = 'h35f7;
        exp_im_rom[605] = 'h7ff66a9;
        exp_im_rom[606] = 'h7fa8c6a;
        exp_im_rom[607] = 'h5470c;
        exp_im_rom[608] = 'h331f0;
        exp_im_rom[609] = 'h3798a;
        exp_im_rom[610] = 'h8ccdc;
        exp_im_rom[611] = 'h7fbed4f;
        exp_im_rom[612] = 'h7fec687;
        exp_im_rom[613] = 'h7ff4a2c;
        exp_im_rom[614] = 'h7fee664;
        exp_im_rom[615] = 'h88b5;
        exp_im_rom[616] = 'h4109;
        exp_im_rom[617] = 'h46a4;
        exp_im_rom[618] = 'ha620;
        exp_im_rom[619] = 'h7ffbfa9;
        exp_im_rom[620] = 'h857;
        exp_im_rom[621] = 'h3739;
        exp_im_rom[622] = 'h108ac;
        exp_im_rom[623] = 'h7ff0511;
        exp_im_rom[624] = 'h7ff99d0;
        exp_im_rom[625] = 'h7ffcd57;
        exp_im_rom[626] = 'h57e3;
        exp_im_rom[627] = 'h7ff1dad;
        exp_im_rom[628] = 'h7ff99a1;
        exp_im_rom[629] = 'hc45;
        exp_im_rom[630] = 'h295b0;
        exp_im_rom[631] = 'h7faf737;
        exp_im_rom[632] = 'h7fcb3c2;
        exp_im_rom[633] = 'h7fc24f7;
        exp_im_rom[634] = 'h7f79263;
        exp_im_rom[635] = 'h444c4;
        exp_im_rom[636] = 'h7ffa77b;
        exp_im_rom[637] = 'h7fd6505;
        exp_im_rom[638] = 'h7f58c79;
        exp_im_rom[639] = 'hbdeac;
        exp_im_rom[640] = 'h4ac7d;
        exp_im_rom[641] = 'h3d7c6;
        exp_im_rom[642] = 'h763cb;
        exp_im_rom[643] = 'h7f89ac0;
        exp_im_rom[644] = 'h7fc41c8;
        exp_im_rom[645] = 'h7faf556;
        exp_im_rom[646] = 'h7f0f329;
        exp_im_rom[647] = 'h12ee9e;
        exp_im_rom[648] = 'h78688;
        exp_im_rom[649] = 'h66f8f;
        exp_im_rom[650] = 'hb0817;
        exp_im_rom[651] = 'h7f7dd2d;
        exp_im_rom[652] = 'h7fe8261;
        exp_im_rom[653] = 'h7ffc811;
        exp_im_rom[654] = 'h16efe;
        exp_im_rom[655] = 'h7fc88a6;
        exp_im_rom[656] = 'h7fe41c1;
        exp_im_rom[657] = 'h7fe24cf;
        exp_im_rom[658] = 'h7fc58cd;
        exp_im_rom[659] = 'h312d4;
        exp_im_rom[660] = 'h2925;
        exp_im_rom[661] = 'h7ff455f;
        exp_im_rom[662] = 'h7fd917d;
        exp_im_rom[663] = 'h24ce2;
        exp_im_rom[664] = 'h7ff9c25;
        exp_im_rom[665] = 'h7fe288e;
        exp_im_rom[666] = 'h7f9ccd1;
        exp_im_rom[667] = 'h99da0;
        exp_im_rom[668] = 'h203ba;
        exp_im_rom[669] = 'h7ff977a;
        exp_im_rom[670] = 'h7f9bed9;
        exp_im_rom[671] = 'h10bef2;
        exp_im_rom[672] = 'h673cf;
        exp_im_rom[673] = 'h548c5;
        exp_im_rom[674] = 'h7249d;
        exp_im_rom[675] = 'h7faa8f6;
        exp_im_rom[676] = 'h7ffcdc3;
        exp_im_rom[677] = 'h1920;
        exp_im_rom[678] = 'h7fe9de9;
        exp_im_rom[679] = 'h75572;
        exp_im_rom[680] = 'h39480;
        exp_im_rom[681] = 'h3a821;
        exp_im_rom[682] = 'h61cb8;
        exp_im_rom[683] = 'h7f88501;
        exp_im_rom[684] = 'h7ff3193;
        exp_im_rom[685] = 'h2848;
        exp_im_rom[686] = 'hbe29;
        exp_im_rom[687] = 'h7ffac9f;
        exp_im_rom[688] = 'h7859;
        exp_im_rom[689] = 'hba83;
        exp_im_rom[690] = 'h13be0;
        exp_im_rom[691] = 'h7fedf18;
        exp_im_rom[692] = 'h371a;
        exp_im_rom[693] = 'h778c;
        exp_im_rom[694] = 'hdcb1;
        exp_im_rom[695] = 'h7fe9ed2;
        exp_im_rom[696] = 'h7ffb4c3;
        exp_im_rom[697] = 'h7ff8099;
        exp_im_rom[698] = 'h7fe182f;
        exp_im_rom[699] = 'h7d68a;
        exp_im_rom[700] = 'h2589b;
        exp_im_rom[701] = 'h1b3ca;
        exp_im_rom[702] = 'h13396;
        exp_im_rom[703] = 'h42539;
        exp_im_rom[704] = 'h2cb6b;
        exp_im_rom[705] = 'h36b67;
        exp_im_rom[706] = 'h673f7;
        exp_im_rom[707] = 'h7ef2d74;
        exp_im_rom[708] = 'h7fd5187;
        exp_im_rom[709] = 'h7fea962;
        exp_im_rom[710] = 'h7fe90c3;
        exp_im_rom[711] = 'h4d9d6;
        exp_im_rom[712] = 'h18304;
        exp_im_rom[713] = 'h1af8b;
        exp_im_rom[714] = 'h31572;
        exp_im_rom[715] = 'h7f6f0e7;
        exp_im_rom[716] = 'h7ff0d5b;
        exp_im_rom[717] = 'ha89;
        exp_im_rom[718] = 'h11b8e;
        exp_im_rom[719] = 'h7fa2836;
        exp_im_rom[720] = 'h7ff2293;
        exp_im_rom[721] = 'h7ffb7a2;
        exp_im_rom[722] = 'h3701;
        exp_im_rom[723] = 'h7fd8e91;
        exp_im_rom[724] = 'h7ffa61c;
        exp_im_rom[725] = 'h7fff6b0;
        exp_im_rom[726] = 'h62e6;
        exp_im_rom[727] = 'h7fcec13;
        exp_im_rom[728] = 'h7ff8f7b;
        exp_im_rom[729] = 'h7ffd970;
        exp_im_rom[730] = 'h29d1;
        exp_im_rom[731] = 'h7fd739d;
        exp_im_rom[732] = 'h7ff920f;
        exp_im_rom[733] = 'h7ffc538;
        exp_im_rom[734] = 'h7fffc17;
        exp_im_rom[735] = 'h7fd8e21;
        exp_im_rom[736] = 'h7ff64e5;
        exp_im_rom[737] = 'h7ff6723;
        exp_im_rom[738] = 'h7ff1434;
        exp_im_rom[739] = 'h4eab7;
        exp_im_rom[740] = 'h343c;
        exp_im_rom[741] = 'h7ffcc9b;
        exp_im_rom[742] = 'h7ff28ae;
        exp_im_rom[743] = 'ha2386;
        exp_im_rom[744] = 'h112ab;
        exp_im_rom[745] = 'ha12d;
        exp_im_rom[746] = 'h6c57;
        exp_im_rom[747] = 'h1cbce;
        exp_im_rom[748] = 'h8d59;
        exp_im_rom[749] = 'h83f5;
        exp_im_rom[750] = 'h9aad;
        exp_im_rom[751] = 'h7fcffc3;
        exp_im_rom[752] = 'h1ff8;
        exp_im_rom[753] = 'h3888;
        exp_im_rom[754] = 'h4180;
        exp_im_rom[755] = 'h549c;
        exp_im_rom[756] = 'h505b;
        exp_im_rom[757] = 'h5bc1;
        exp_im_rom[758] = 'h7a8e;
        exp_im_rom[759] = 'h7fa82f4;
        exp_im_rom[760] = 'h1e35;
        exp_im_rom[761] = 'h45b3;
        exp_im_rom[762] = 'h794f;
        exp_im_rom[763] = 'h7f01072;
        exp_im_rom[764] = 'h7ffe4e2;
        exp_im_rom[765] = 'h15e9;
        exp_im_rom[766] = 'h3b31;
        exp_im_rom[767] = 'h7d74a2a;
        exp_im_rom[768] = 'h10;
        exp_im_rom[769] = 'h267f;
        exp_im_rom[770] = 'h5d1a;
        exp_im_rom[771] = 'h1e9dd0;
        exp_im_rom[772] = 'h7ffb427;
        exp_im_rom[773] = 'h7fff3c0;
        exp_im_rom[774] = 'h3a6d;
        exp_im_rom[775] = 'h121401;
        exp_im_rom[776] = 'h7ff2cb3;
        exp_im_rom[777] = 'h7ff5bf2;
        exp_im_rom[778] = 'h7ff4258;
        exp_im_rom[779] = 'h7f92161;
        exp_im_rom[780] = 'h7ffa07a;
        exp_im_rom[781] = 'h7ff2fbf;
        exp_im_rom[782] = 'h7fe41c8;
        exp_im_rom[783] = 'h7df3954;
        exp_im_rom[784] = 'h21394;
        exp_im_rom[785] = 'hfaa8;
        exp_im_rom[786] = 'h8def;
        exp_im_rom[787] = 'h7fe9892;
        exp_im_rom[788] = 'h7cbc;
        exp_im_rom[789] = 'h3f64;
        exp_im_rom[790] = 'h7ffecf4;
        exp_im_rom[791] = 'h7fa79d3;
        exp_im_rom[792] = 'hd6f0;
        exp_im_rom[793] = 'h6e44;
        exp_im_rom[794] = 'h1e28;
        exp_im_rom[795] = 'h7fc9c43;
        exp_im_rom[796] = 'hb3ec;
        exp_im_rom[797] = 'h4850;
        exp_im_rom[798] = 'h7ffb93a;
        exp_im_rom[799] = 'h7f70f74;
        exp_im_rom[800] = 'h228fd;
        exp_im_rom[801] = 'h19422;
        exp_im_rom[802] = 'h1ca04;
        exp_im_rom[803] = 'h8c002;
        exp_im_rom[804] = 'h7ff520a;
        exp_im_rom[805] = 'h7fff381;
        exp_im_rom[806] = 'h2161;
        exp_im_rom[807] = 'ha963;
        exp_im_rom[808] = 'h7fff7c5;
        exp_im_rom[809] = 'h7fff2e8;
        exp_im_rom[810] = 'h7ffbe7e;
        exp_im_rom[811] = 'h7fd0613;
        exp_im_rom[812] = 'hcb33;
        exp_im_rom[813] = 'h61f2;
        exp_im_rom[814] = 'h2626;
        exp_im_rom[815] = 'h7ff01db;
        exp_im_rom[816] = 'h59fc;
        exp_im_rom[817] = 'h7fff782;
        exp_im_rom[818] = 'h7ff59b8;
        exp_im_rom[819] = 'h7f95b7e;
        exp_im_rom[820] = 'h22d4c;
        exp_im_rom[821] = 'h11152;
        exp_im_rom[822] = 'h7f4c;
        exp_im_rom[823] = 'h7fd9f70;
        exp_im_rom[824] = 'h1afa8;
        exp_im_rom[825] = 'h10677;
        exp_im_rom[826] = 'h95e9;
        exp_im_rom[827] = 'h7fe2efd;
        exp_im_rom[828] = 'h19e0f;
        exp_im_rom[829] = 'hd2cc;
        exp_im_rom[830] = 'h7ffc458;
        exp_im_rom[831] = 'h7f62d36;
        exp_im_rom[832] = 'h6b17b;
        exp_im_rom[833] = 'h51d4b;
        exp_im_rom[834] = 'h65039;
        exp_im_rom[835] = 'h1584da;
        exp_im_rom[836] = 'h7fb0152;
        exp_im_rom[837] = 'h7ff147a;
        exp_im_rom[838] = 'h871a;
        exp_im_rom[839] = 'h45928;
        exp_im_rom[840] = 'h7fed300;
        exp_im_rom[841] = 'h18ce;
        exp_im_rom[842] = 'hd306;
        exp_im_rom[843] = 'h366d2;
        exp_im_rom[844] = 'h7ff939f;
        exp_im_rom[845] = 'hc0bd;
        exp_im_rom[846] = 'h1eebe;
        exp_im_rom[847] = 'h8c7ed;
        exp_im_rom[848] = 'h7fc6089;
        exp_im_rom[849] = 'h7ff03cf;
        exp_im_rom[850] = 'h6674;
        exp_im_rom[851] = 'h69a41;
        exp_im_rom[852] = 'h7fab1f1;
        exp_im_rom[853] = 'h7fcb53c;
        exp_im_rom[854] = 'h7fc580f;
        exp_im_rom[855] = 'h7f595af;
        exp_im_rom[856] = 'h43f17;
        exp_im_rom[857] = 'h176ab;
        exp_im_rom[858] = 'h103bd;
        exp_im_rom[859] = 'h26d23;
        exp_im_rom[860] = 'h7fe48c9;
        exp_im_rom[861] = 'h7fea11c;
        exp_im_rom[862] = 'h7fdc778;
        exp_im_rom[863] = 'h7f77461;
        exp_im_rom[864] = 'h55fe9;
        exp_im_rom[865] = 'h21ae9;
        exp_im_rom[866] = 'h10ffa;
        exp_im_rom[867] = 'h7feab93;
        exp_im_rom[868] = 'h3680f;
        exp_im_rom[869] = 'h24886;
        exp_im_rom[870] = 'h24867;
        exp_im_rom[871] = 'h416d1;
        exp_im_rom[872] = 'h7ff63a9;
        exp_im_rom[873] = 'h84c7;
        exp_im_rom[874] = 'hcb6b;
        exp_im_rom[875] = 'h1241b;
        exp_im_rom[876] = 'h97e1;
        exp_im_rom[877] = 'hcc3b;
        exp_im_rom[878] = 'hdfcd;
        exp_im_rom[879] = 'hf0a6;
        exp_im_rom[880] = 'hfc44;
        exp_im_rom[881] = 'h1170f;
        exp_im_rom[882] = 'h154f2;
        exp_im_rom[883] = 'h2d50a;
        exp_im_rom[884] = 'h7fe5dc8;
        exp_im_rom[885] = 'h7ff23f3;
        exp_im_rom[886] = 'h7fe24f2;
        exp_im_rom[887] = 'h7f6ddd5;
        exp_im_rom[888] = 'hc306e;
        exp_im_rom[889] = 'h6486b;
        exp_im_rom[890] = 'h5b185;
        exp_im_rom[891] = 'h76898;
        exp_im_rom[892] = 'h31750;
        exp_im_rom[893] = 'h6118f;
        exp_im_rom[894] = 'ha129b;
        exp_im_rom[895] = 'h1d9234;
        exp_im_rom[896] = 'h7e2cc71;
        exp_im_rom[897] = 'h7f5ab8e;
        exp_im_rom[898] = 'h7f83909;
        exp_im_rom[899] = 'h7f2e375;
        exp_im_rom[900] = 'ha6455;
        exp_im_rom[901] = 'h3aaf8;
        exp_im_rom[902] = 'h3670d;
        exp_im_rom[903] = 'h6a15e;
        exp_im_rom[904] = 'h7fbad17;
        exp_im_rom[905] = 'h7fffe07;
        exp_im_rom[906] = 'h17c7d;
        exp_im_rom[907] = 'h4b698;
        exp_im_rom[908] = 'h7fc52a4;
        exp_im_rom[909] = 'h84d4;
        exp_im_rom[910] = 'h2d4fc;
        exp_im_rom[911] = 'ha70e6;
        exp_im_rom[912] = 'h7f0bbc7;
        exp_im_rom[913] = 'h7fadcae;
        exp_im_rom[914] = 'h7fc7aae;
        exp_im_rom[915] = 'h7fb9a0c;
        exp_im_rom[916] = 'h34d81;
        exp_im_rom[917] = 'h12b90;
        exp_im_rom[918] = 'h1af2e;
        exp_im_rom[919] = 'h4c52f;
        exp_im_rom[920] = 'h7f95684;
        exp_im_rom[921] = 'h7fe9953;
        exp_im_rom[922] = 'h214d;
        exp_im_rom[923] = 'h3123c;
        exp_im_rom[924] = 'h7f98dac;
        exp_im_rom[925] = 'h7fe672d;
        exp_im_rom[926] = 'h2e0;
        exp_im_rom[927] = 'h3ad14;
        exp_im_rom[928] = 'h7f5bc98;
        exp_im_rom[929] = 'h7fc4952;
        exp_im_rom[930] = 'h7fd552f;
        exp_im_rom[931] = 'h7fd5819;
        exp_im_rom[932] = 'h51c7;
        exp_im_rom[933] = 'h7ff7fad;
        exp_im_rom[934] = 'h7ffdda4;
        exp_im_rom[935] = 'h18972;
        exp_im_rom[936] = 'h7f9bdf9;
        exp_im_rom[937] = 'h7fd95b2;
        exp_im_rom[938] = 'h7fe20f7;
        exp_im_rom[939] = 'h7fe1b15;
        exp_im_rom[940] = 'h7ffd46e;
        exp_im_rom[941] = 'h7ff2e78;
        exp_im_rom[942] = 'h7ff2fb7;
        exp_im_rom[943] = 'h7ff49d4;
        exp_im_rom[944] = 'h7ff0983;
        exp_im_rom[945] = 'h7ff46eb;
        exp_im_rom[946] = 'h7ff6bc9;
        exp_im_rom[947] = 'h7ffcf4c;
        exp_im_rom[948] = 'h7fdb7e2;
        exp_im_rom[949] = 'h7fec735;
        exp_im_rom[950] = 'h7fea9b6;
        exp_im_rom[951] = 'h7fd549a;
        exp_im_rom[952] = 'h7898c;
        exp_im_rom[953] = 'h2a329;
        exp_im_rom[954] = 'h339b3;
        exp_im_rom[955] = 'h7a556;
        exp_im_rom[956] = 'h7e92908;
        exp_im_rom[957] = 'h7fab529;
        exp_im_rom[958] = 'h7fce310;
        exp_im_rom[959] = 'h7fe8219;
        exp_im_rom[960] = 'h7f78e06;
        exp_im_rom[961] = 'h7fba0cc;
        exp_im_rom[962] = 'h7fb619f;
        exp_im_rom[963] = 'h7f88e24;
        exp_im_rom[964] = 'hfc7f1;
        exp_im_rom[965] = 'h18182;
        exp_im_rom[966] = 'h7ffea7d;
        exp_im_rom[967] = 'h7fee84f;
        exp_im_rom[968] = 'h1df1d;
        exp_im_rom[969] = 'h7ff53fe;
        exp_im_rom[970] = 'h7fe7975;
        exp_im_rom[971] = 'h7fc5beb;
        exp_im_rom[972] = 'hde2f9;
        exp_im_rom[973] = 'h242d2;
        exp_im_rom[974] = 'h1469a;
        exp_im_rom[975] = 'h15a3e;
        exp_im_rom[976] = 'h7fbaec3;
        exp_im_rom[977] = 'h7ff11e0;
        exp_im_rom[978] = 'h7ff0380;
        exp_im_rom[979] = 'h7fe26de;
        exp_im_rom[980] = 'h78e83;
        exp_im_rom[981] = 'hda6d;
        exp_im_rom[982] = 'h3894;
        exp_im_rom[983] = 'h7ffb715;
        exp_im_rom[984] = 'h2d3c5;
        exp_im_rom[985] = 'h4b29;
        exp_im_rom[986] = 'h7ffdec8;
        exp_im_rom[987] = 'h7ff049d;
        exp_im_rom[988] = 'h9bdac;
        exp_im_rom[989] = 'h1cbdc;
        exp_im_rom[990] = 'h1883d;
        exp_im_rom[991] = 'h248d4;
        exp_im_rom[992] = 'h7f3cf3e;
        exp_im_rom[993] = 'h7fee892;
        exp_im_rom[994] = 'h7ff89be;
        exp_im_rom[995] = 'h7ffcd82;
        exp_im_rom[996] = 'h7fedee3;
        exp_im_rom[997] = 'h7ffc4c4;
        exp_im_rom[998] = 'h7ffe0e7;
        exp_im_rom[999] = 'h79f;
        exp_im_rom[1000] = 'h7fdb2f1;
        exp_im_rom[1001] = 'h7ffa955;
        exp_im_rom[1002] = 'h7ffc2b4;
        exp_im_rom[1003] = 'h7ffcd51;
        exp_im_rom[1004] = 'h7ffc2f6;
        exp_im_rom[1005] = 'h7ffd456;
        exp_im_rom[1006] = 'h7ffd787;
        exp_im_rom[1007] = 'h7ffd9d7;
        exp_im_rom[1008] = 'h7ffd163;
        exp_im_rom[1009] = 'h7ffdab4;
        exp_im_rom[1010] = 'h7ffdab3;
        exp_im_rom[1011] = 'h7ffd74a;
        exp_im_rom[1012] = 'h8acb;
        exp_im_rom[1013] = 'h7ffe77d;
        exp_im_rom[1014] = 'h7ffe19f;
        exp_im_rom[1015] = 'h7ffd749;
        exp_im_rom[1016] = 'h25b76;
        exp_im_rom[1017] = 'h7ffff50;
        exp_im_rom[1018] = 'h7fff5f3;
        exp_im_rom[1019] = 'h7fff083;
        exp_im_rom[1020] = 'h1cd55;
        exp_im_rom[1021] = 'h16;
        exp_im_rom[1022] = 'h7fffdbd;
        exp_im_rom[1023] = 'h7fffe42;
    end
end
initial begin
    fft_blk_exp[0] = 'h0;
    ifft_blk_exp[0] = 'h0;
end



always @(posedge i_clk or negedge i_rstn) begin
    if (~i_rstn) begin
        o_rdata <= {(OUTPUT_WIDTH*2){1'b0}};
    end        
    else if (i_clken) begin
        o_rdata[OUTPUT_WIDTH-1:0] <= exp_re_rom[i_addr];
        o_rdata[OUTPUT_WIDTH*2-1:OUTPUT_WIDTH] <= exp_im_rom[i_addr];
    end
end
      
assign o_blk_exp = FFT_MODE ? fft_blk_exp[0] : ifft_blk_exp[0];

endmodule