module x(
        input wire [10:0]i,
        output reg [15:0] data
   );
always @(*) begin
case(i)
   0 :   data= -180 ;
   1 :   data= -116 ;
   2 :   data= -136 ;
   3 :   data= -155 ;
   4 :   data= -174 ;
   5 :   data= -212 ;
   6 :   data= -192 ;
   7 :   data= -96 ;
   8 :   data= -57 ;
   9 :   data= -109 ;
   10 :  data= -127 ;
   11 :  data= -75 ;
   12 :  data= -13 ;
   13 :  data= 73 ;
   14 :  data= 163 ;
   15 :  data= 166 ;
   16 :  data= 127 ;
   17 :  data= 156 ;
   18 :  data= 202 ;
   19 :  data= 196 ;
   20 :  data= 195 ;
   21 :  data= 221 ;
   22 :  data= 234 ;
   23 :  data= 238 ;
   24 :  data= 245 ;
   25 :  data= 250 ;
   26 :  data= 276 ;
   27 :  data= 283 ;
   28 :  data= 215 ;
   29 :  data= 153 ;
   30 :  data= 157 ;
   31 :  data= 115 ;
   32 :  data= -7 ;
   33 :  data= -61 ;
   34 :  data= -30 ;
   35 :  data= -73 ;
   36 :  data= -180 ;
   37 :  data= -191 ;
   38 :  data= -114 ;
   39 :  data= -96 ;
   40 :  data= -162 ;
   41 :  data= -212 ;
   42 :  data= -181 ;
   43 :  data= -115 ;
   44 :  data= -103 ;
   45 :  data= -129 ;
   46 :  data= -91 ;
   47 :  data= 14 ;
   48 :  data= 75 ;
   49 :  data= 32 ;
   50 :  data= -88 ;
   51 :  data= -223 ;
   52 :  data= -267 ;
   53 :  data= -204 ;
   54 :  data= -156 ;
   55 :  data= -169 ;
   56 :  data= -168 ;
   57 :  data= -148 ;
   58 :  data= -147 ;
   59 :  data= -118 ;
   60 :  data= -53 ;
   61 :  data= -22 ;
   62 :  data= -29 ;
   63 :  data= -30 ;
   64 :  data= -26 ;
   65 :  data= -18 ;
   66 :  data= -12 ;
   67 :  data= -49 ;
   68 :  data= -110 ;
   69 :  data= -120 ;
   70 :  data= -107 ;
   71 :  data= -149 ;
   72 :  data= -228 ;
   73 :  data= -260 ;
   74 :  data= -217 ;
   75 :  data= -160 ;
   76 :  data= -180 ;
   77 :  data= -261 ;
   78 :  data= -304 ;
   79 :  data= -301 ;
   80 :  data= -298 ;
   81 :  data= -250 ;
   82 :  data= -149 ;
   83 :  data= -120 ;
   84 :  data= -207 ;
   85 :  data= -301 ;
   86 :  data= -352 ;
   87 :  data= -398 ;
   88 :  data= -435 ;
   89 :  data= -460 ;
   90 :  data= -488 ;
   91 :  data= -495 ;
   92 :  data= -458 ;
   93 :  data= -410 ;
   94 :  data= -399 ;
   95 :  data= -444 ;
   96 :  data= -513 ;
   97 :  data= -534 ;
   98 :  data= -509 ;
   99 :  data= -500 ;
   100 :  data=-501 ;
   101 :  data=-479 ;
   102 :  data=-453 ;
   103 :  data=-392 ;
   104 :  data=-274 ;
   105 :  data=-207 ;
   106 :  data=-210 ;
   107 :  data=-114 ;
   108 :  data=96 ;
   109 :  data=214 ;
   110 :  data=189 ;
   111 :  data=167 ;
   112 :  data=200 ;
   113 :  data=214 ;
   114 :  data=187 ;
   115 :  data=190 ;
   116 :  data=272 ;
   117 :  data=335 ;
   118 :  data=274 ;
   119 :  data=183 ;
   120 :  data=174 ;
   121 :  data=151 ;
   122 :  data=62 ;
   123 :  data=40 ;
   124 :  data=78 ;
   125 :  data=33 ;
   126 :  data=-34 ;
   127 :  data=6 ;
   128 :  data=66 ;
   129 :  data=35 ;
   130 :  data=-6 ;
   131 :  data=27 ;
   132 :  data=111 ;
   133 :  data=173 ;
   134 :  data=150 ;
   135 :  data=76 ;
   136 :  data=39 ;
   137 :  data=4 ;
   138 :  data=-91 ;
   139 :  data=-136 ;
   140 :  data=-69 ;
   141 :  data=-59 ;
   142 :  data=-148 ;
   143 :  data=-149 ;
   144 :  data=-71 ;
   145 :  data=-104 ;
   146 :  data=-201 ;
   147 :  data=-193 ;
   148 :  data=-130 ;
   149 :  data=-101 ;
   150 :  data=-44 ;
   151 :  data=28 ;
   152 :  data=19 ;
   153 :  data=-16 ;
   154 :  data=21 ;
   155 :  data=75 ;
   156 :  data=84 ;
   157 :  data=94 ;
   158 :  data=111 ;
   159 :  data=105 ;
   160 :  data=129 ;
   161 :  data=199 ;
   162 :  data=219 ;
   163 :  data=158 ;
   164 :  data=109 ;
   165 :  data=129 ;
   166 :  data=183 ;
   167 :  data=216 ;
   168 :  data=197 ;
   169 :  data=148 ;
   170 :  data=125 ;
   171 :  data=136 ;
   172 :  data=146 ;
   173 :  data=163 ;
   174 :  data=225 ;
   175 :  data=291 ;
   176 :  data=279 ;
   177 :  data=232 ;
   178 :  data=251 ;
   179 :  data=304 ;
   180 :  data=295 ;
   181 :  data=250 ;
   182 :  data=238 ;
   183 :  data=242 ;
   184 :  data=243 ;
   185 :  data=245 ;
   186 :  data=206 ;
   187 :  data=134 ;
   188 :  data=136 ;
   189 :  data=224 ;
   190 :  data=286 ;
   191 :  data=289 ;
   192 :  data=282 ;
   193 :  data=267 ;
   194 :  data=259 ;
   195 :  data=307 ;
   196 :  data=366 ;
   197 :  data=353 ;
   198 :  data=293 ;
   199 :  data=266 ;
   200 :  data=279 ;
   201 :  data=283 ;
   202 :  data=241 ;
   203 :  data=173 ;
   204 :  data=136 ;
   205 :  data=138 ;
   206 :  data=161 ;
   207 :  data=213 ;
   208 :  data=258 ;
   209 :  data=223 ;
   210 :  data=153 ;
   211 :  data=163 ;
   212 :  data=219 ;
   213 :  data=224 ;
   214 :  data=221 ;
   215 :  data=258 ;
   216 :  data=272 ;
   217 :  data=262 ;
   218 :  data=326 ;
   219 :  data=442 ;
   220 :  data=484 ;
   221 :  data=438 ;
   222 :  data=399 ;
   223 :  data=412 ;
   224 :  data=466 ;
   225 :  data=530 ;
   226 :  data=539 ;
   227 :  data=465 ;
   228 :  data=394 ;
   229 :  data=421 ;
   230 :  data=498 ;
   231 :  data=507 ;
   232 :  data=464 ;
   233 :  data=486 ;
   234 :  data=560 ;
   235 :  data=561 ;
   236 :  data=520 ;
   237 :  data=564 ;
   238 :  data=620 ;
   239 :  data=572 ;
   240 :  data=548 ;
   241 :  data=641 ;
   242 :  data=667 ;
   243 :  data=537 ;
   244 :  data=439 ;
   245 :  data=447 ;
   246 :  data=439 ;
   247 :  data=402 ;
   248 :  data=395 ;
   249 :  data=373 ;
   250 :  data=326 ;
   251 :  data=309 ;
   252 :  data=308 ;
   253 :  data=298 ;
   254 :  data=315 ;
   255 :  data=358 ;
   256 :  data=388 ;
   257 :  data=411 ;
   258 :  data=436 ;
   259 :  data=465 ;
   260 :  data=512 ;
   261 :  data=559 ;
   262 :  data=579 ;
   263 :  data=603 ;
   264 :  data=644 ;
   265 :  data=641 ;
   266 :  data=586 ;
   267 :  data=558 ;
   268 :  data=577 ;
   269 :  data=574 ;
   270 :  data=526 ;
   271 :  data=509 ;
   272 :  data=564 ;
   273 :  data=591 ;
   274 :  data=521 ;
   275 :  data=455 ;
   276 :  data=466 ;
   277 :  data=474 ;
   278 :  data=461 ;
   279 :  data=508 ;
   280 :  data=571 ;
   281 :  data=567 ;
   282 :  data=555 ;
   283 :  data=574 ;
   284 :  data=570 ;
   285 :  data=576 ;
   286 :  data=631 ;
   287 :  data=618 ;
   288 :  data=492 ;
   289 :  data=425 ;
   290 :  data=498 ;
   291 :  data=542 ;
   292 :  data=450 ;
   293 :  data=350 ;
   294 :  data=349 ;
   295 :  data=370 ;
   296 :  data=356 ;
   297 :  data=375 ;
   298 :  data=428 ;
   299 :  data=412 ;
   300 :  data=322 ;
   301 :  data=252 ;
   302 :  data=248 ;
   303 :  data=328 ;
   304 :  data=490 ;
   305 :  data=618 ;
   306 :  data=626 ;
   307 :  data=610 ;
   308 :  data=639 ;
   309 :  data=636 ;
   310 :  data=604 ;
   311 :  data=644 ;
   312 :  data=723 ;
   313 :  data=712 ;
   314 :  data=638 ;
   315 :  data=629 ;
   316 :  data=698 ;
   317 :  data=761 ;
   318 :  data=806 ;
   319 :  data=907 ;
   320 :  data=1066 ;
   321 :  data=1166 ;
   322 :  data=1150 ;
   323 :  data=1115 ;
   324 :  data=1154 ;
   325 :  data=1210 ;
   326 :  data=1210 ;
   327 :  data=1188 ;
   328 :  data=1162 ;
   329 :  data=1053 ;
   330 :  data=897 ;
   331 :  data=880 ;
   332 :  data=1009 ;
   333 :  data=1075 ;
   334 :  data=1024 ;
   335 :  data=989 ;
   336 :  data=993 ;
   337 :  data=971 ;
   338 :  data=943 ;
   339 :  data=933 ;
   340 :  data=923 ;
   341 :  data=922 ;
   342 :  data=911 ;
   343 :  data=856 ;
   344 :  data=806 ;
   345 :  data=794 ;
   346 :  data=767 ;
   347 :  data=734 ;
   348 :  data=742 ;
   349 :  data=766 ;
   350 :  data=800 ;
   351 :  data=842 ;
   352 :  data=801 ;
   353 :  data=689 ;
   354 :  data=665 ;
   355 :  data=713 ;
   356 :  data=673 ;
   357 :  data=572 ;
   358 :  data=535 ;
   359 :  data=547 ;
   360 :  data=557 ;
   361 :  data=543 ;
   362 :  data=470 ;
   363 :  data=388 ;
   364 :  data=383 ;
   365 :  data=410 ;
   366 :  data=401 ;
   367 :  data=389 ;
   368 :  data=396 ;
   369 :  data=383 ;
   370 :  data=360 ;
   371 :  data=374 ;
   372 :  data=444 ;
   373 :  data=540 ;
   374 :  data=600 ;
   375 :  data=606 ;
   376 :  data=597 ;
   377 :  data=592 ;
   378 :  data=579 ;
   379 :  data=564 ;
   380 :  data=537 ;
   381 :  data=518 ;
   382 :  data=556 ;
   383 :  data=593 ;
   384 :  data=537 ;
   385 :  data=445 ;
   386 :  data=400 ;
   387 :  data=375 ;
   388 :  data=376 ;
   389 :  data=425 ;
   390 :  data=444 ;
   391 :  data=426 ;
   392 :  data=450 ;
   393 :  data=459 ;
   394 :  data=392 ;
   395 :  data=363 ;
   396 :  data=414 ;
   397 :  data=446 ;
   398 :  data=460 ;
   399 :  data=496 ;
   400 :  data=500 ;
   401 :  data=486 ;
   402 :  data=519 ;
   403 :  data=549 ;
   404 :  data=542 ;
   405 :  data=552 ;
   406 :  data=564 ;
   407 :  data=549 ;
   408 :  data=557 ;
   409 :  data=554 ;
   410 :  data=452 ;
   411 :  data=348 ;
   412 :  data=373 ;
   413 :  data=439 ;
   414 :  data=458 ;
   415 :  data=477 ;
   416 :  data=474 ;
   417 :  data=394 ;
   418 :  data=349 ;
   419 :  data=443 ;
   420 :  data=573 ;
   421 :  data=673 ;
   422 :  data=810 ;
   423 :  data=931 ;
   424 :  data=922 ;
   425 :  data=881 ;
   426 :  data=920 ;
   427 :  data=940 ;
   428 :  data=888 ;
   429 :  data=874 ;
   430 :  data=888 ;
   431 :  data=816 ;
   432 :  data=707 ;
   433 :  data=667 ;
   434 :  data=669 ;
   435 :  data=663 ;
   436 :  data=649 ;
   437 :  data=626 ;
   438 :  data=612 ;
   439 :  data=614 ;
   440 :  data=587 ;
   441 :  data=528 ;
   442 :  data=475 ;
   443 :  data=406 ;
   444 :  data=334 ;
   445 :  data=334 ;
   446 :  data=370 ;
   447 :  data=359 ;
   448 :  data=335 ;
   449 :  data=326 ;
   450 :  data=269 ;
   451 :  data=171 ;
   452 :  data=123 ;
   453 :  data=132 ;
   454 :  data=163 ;
   455 :  data=226 ;
   456 :  data=308 ;
   457 :  data=331 ;
   458 :  data=254 ;
   459 :  data=166 ;
   460 :  data=170 ;
   461 :  data=233 ;
   462 :  data=265 ;
   463 :  data=296 ;
   464 :  data=355 ;
   465 :  data=379 ;
   466 :  data=372 ;
   467 :  data=397 ;
   468 :  data=415 ;
   469 :  data=397 ;
   470 :  data=399 ;
   471 :  data=386 ;
   472 :  data=326 ;
   473 :  data=334 ;
   474 :  data=410 ;
   475 :  data=413 ;
   476 :  data=394 ;
   477 :  data=434 ;
   478 :  data=377 ;
   479 :  data=191 ;
   480 :  data=112 ;
   481 :  data=145 ;
   482 :  data=94 ;
   483 :  data=9 ;
   484 :  data=27 ;
   485 :  data=51 ;
   486 :  data=1 ;
   487 :  data=-45 ;
   488 :  data=-79 ;
   489 :  data=-122 ;
   490 :  data=-90 ;
   491 :  data=43 ;
   492 :  data=178 ;
   493 :  data=275 ;
   494 :  data=343 ;
   495 :  data=313 ;
   496 :  data=165 ;
   497 :  data=54 ;
   498 :  data=72 ;
   499 :  data=105 ;
   500 :  data=76 ;
   501 :  data=60 ;
   502 :  data=39 ;
   503 :  data=-101 ;
   504 :  data=-304 ;
   505 :  data=-427 ;
   506 :  data=-504 ;
   507 :  data=-582 ;
   508 :  data=-557 ;
   509 :  data=-442 ;
   510 :  data=-409 ;
   511 :  data=-446 ;
   512 :  data=-416 ;
   513 :  data=-365 ;
   514 :  data=-363 ;
   515 :  data=-316 ;
   516 :  data=-231 ;
   517 :  data=-241 ;
   518 :  data=-290 ;
   519 :  data=-247 ;
   520 :  data=-212 ;
   521 :  data=-279 ;
   522 :  data=-310 ;
   523 :  data=-238 ;
   524 :  data=-202 ;
   525 :  data=-253 ;
   526 :  data=-300 ;
   527 :  data=-316 ;
   528 :  data=-336 ;
   529 :  data=-362 ;
   530 :  data=-392 ;
   531 :  data=-413 ;
   532 :  data=-402 ;
   533 :  data=-370 ;
   534 :  data=-320 ;
   535 :  data=-255 ;
   536 :  data=-251 ;
   537 :  data=-355 ;
   538 :  data=-456 ;
   539 :  data=-466 ;
   540 :  data=-455 ;
   541 :  data=-460 ;
   542 :  data=-426 ;
   543 :  data=-377 ;
   544 :  data=-390 ;
   545 :  data=-424 ;
   546 :  data=-410 ;
   547 :  data=-390 ;
   548 :  data=-387 ;
   549 :  data=-298 ;
   550 :  data=-90 ;
   551 :  data=66 ;
   552 :  data=35 ;
   553 :  data=-123 ;
   554 :  data=-312 ;
   555 :  data=-495 ;
   556 :  data=-628 ;
   557 :  data=-683 ;
   558 :  data=-666 ;
   559 :  data=-573 ;
   560 :  data=-485 ;
   561 :  data=-533 ;
   562 :  data=-620 ;
   563 :  data=-572 ;
   564 :  data=-479 ;
   565 :  data=-448 ;
   566 :  data=-354 ;
   567 :  data=-194 ;
   568 :  data=-135 ;
   569 :  data=-141 ;
   570 :  data=-137 ;
   571 :  data=-228 ;
   572 :  data=-375 ;
   573 :  data=-417 ;
   574 :  data=-424 ;
   575 :  data=-474 ;
   576 :  data=-431 ;
   577 :  data=-307 ;
   578 :  data=-265 ;
   579 :  data=-267 ;
   580 :  data=-170 ;
   581 :  data=41 ;
   582 :  data=284 ;
   583 :  data=431 ;
   584 :  data=427 ;
   585 :  data=368 ;
   586 :  data=280 ;
   587 :  data=102 ;
   588 :  data=-59 ;
   589 :  data=-100 ;
   590 :  data=-117 ;
   591 :  data=-121 ;
   592 :  data=-54 ;
   593 :  data=-29 ;
   594 :  data=-61 ;
   595 :  data=0 ;
   596 :  data=70 ;
   597 :  data=7 ;
   598 :  data=-60 ;
   599 :  data=-81 ;
   600 :  data=-151 ;
   601 :  data=-168 ;
   602 :  data=-77 ;
   603 :  data=-87 ;
   604 :  data=-229 ;
   605 :  data=-328 ;
   606 :  data=-374 ;
   607 :  data=-400 ;
   608 :  data=-342 ;
   609 :  data=-233 ;
   610 :  data=-141 ;
   611 :  data=-58 ;
   612 :  data=-37 ;
   613 :  data=-92 ;
   614 :  data=-123 ;
   615 :  data=-166 ;
   616 :  data=-262 ;
   617 :  data=-252 ;
   618 :  data=-85 ;
   619 :  data=88 ;
   620 :  data=226 ;
   621 :  data=303 ;
   622 :  data=228 ;
   623 :  data=94 ;
   624 :  data=44 ;
   625 :  data=34 ;
   626 :  data=89 ;
   627 :  data=275 ;
   628 :  data=410 ;
   629 :  data=409 ;
   630 :  data=456 ;
   631 :  data=549 ;
   632 :  data=546 ;
   633 :  data=555 ;
   634 :  data=649 ;
   635 :  data=673 ;
   636 :  data=624 ;
   637 :  data=603 ;
   638 :  data=526 ;
   639 :  data=367 ;
   640 :  data=268 ;
   641 :  data=235 ;
   642 :  data=187 ;
   643 :  data=166 ;
   644 :  data=203 ;
   645 :  data=232 ;
   646 :  data=237 ;
   647 :  data=261 ;
   648 :  data=318 ;
   649 :  data=362 ;
   650 :  data=309 ;
   651 :  data=149 ;
   652 :  data=2 ;
   653 :  data=-36 ;
   654 :  data=26 ;
   655 :  data=157 ;
   656 :  data=287 ;
   657 :  data=336 ;
   658 :  data=311 ;
   659 :  data=244 ;
   660 :  data=147 ;
   661 :  data=89 ;
   662 :  data=114 ;
   663 :  data=139 ;
   664 :  data=102 ;
   665 :  data=52 ;
   666 :  data=-38 ;
   667 :  data=-256 ;
   668 :  data=-524 ;
   669 :  data=-647 ;
   670 :  data=-564 ;
   671 :  data=-357 ;
   672 :  data=-110 ;
   673 :  data=67 ;
   674 :  data=44 ;
   675 :  data=-133 ;
   676 :  data=-264 ;
   677 :  data=-277 ;
   678 :  data=-243 ;
   679 :  data=-155 ;
   680 :  data=-36 ;
   681 :  data=-33 ;
   682 :  data=-136 ;
   683 :  data=-170 ;
   684 :  data=-150 ;
   685 :  data=-187 ;
   686 :  data=-213 ;
   687 :  data=-215 ;
   688 :  data=-312 ;
   689 :  data=-454 ;
   690 :  data=-506 ;
   691 :  data=-521 ;
   692 :  data=-531 ;
   693 :  data=-447 ;
   694 :  data=-308 ;
   695 :  data=-212 ;
   696 :  data=-138 ;
   697 :  data=-115 ;
   698 :  data=-209 ;
   699 :  data=-301 ;
   700 :  data=-285 ;
   701 :  data=-264 ;
   702 :  data=-272 ;
   703 :  data=-219 ;
   704 :  data=-163 ;
   705 :  data=-222 ;
   706 :  data=-347 ;
   707 :  data=-478 ;
   708 :  data=-608 ;
   709 :  data=-648 ;
   710 :  data=-564 ;
   711 :  data=-488 ;
   712 :  data=-435 ;
   713 :  data=-300 ;
   714 :  data=-230 ;
   715 :  data=-420 ;
   716 :  data=-605 ;
   717 :  data=-442 ;
   718 :  data=-156 ;
   719 :  data=-118 ;
   720 :  data=-171 ;
   721 :  data=-52 ;
   722 :  data=46 ;
   723 :  data=-56 ;
   724 :  data=-123 ;
   725 :  data=1 ;
   726 :  data=133 ;
   727 :  data=203 ;
   728 :  data=318 ;
   729 :  data=392 ;
   730 :  data=313 ;
   731 :  data=240 ;
   732 :  data=290 ;
   733 :  data=332 ;
   734 :  data=335 ;
   735 :  data=390 ;
   736 :  data=419 ;
   737 :  data=338 ;
   738 :  data=288 ;
   739 :  data=339 ;
   740 :  data=355 ;
   741 :  data=262 ;
   742 :  data=71 ;
   743 :  data=-184 ;
   744 :  data=-347 ;
   745 :  data=-297 ;
   746 :  data=-167 ;
   747 :  data=-76 ;
   748 :  data=68 ;
   749 :  data=277 ;
   750 :  data=425 ;
   751 :  data=494 ;
   752 :  data=508 ;
   753 :  data=442 ;
   754 :  data=350 ;
   755 :  data=303 ;
   756 :  data=283 ;
   757 :  data=282 ;
   758 :  data=260 ;
   759 :  data=102 ;
   760 :  data=-126 ;
   761 :  data=-218 ;
   762 :  data=-186 ;
   763 :  data=-160 ;
   764 :  data=-114 ;
   765 :  data=-50 ;
   766 :  data=-67 ;
   767 :  data=-112 ;
   768 :  data=-113 ;
   769 :  data=-184 ;
   770 :  data=-355 ;
   771 :  data=-443 ;
   772 :  data=-377 ;
   773 :  data=-264 ;
   774 :  data=-156 ;
   775 :  data=-30 ;
   776 :  data=82 ;
   777 :  data=152 ;
   778 :  data=215 ;
   779 :  data=288 ;
   780 :  data=310 ;
   781 :  data=237 ;
   782 :  data=150 ;
   783 :  data=155 ;
   784 :  data=214 ;
   785 :  data=217 ;
   786 :  data=150 ;
   787 :  data=80 ;
   788 :  data=44 ;
   789 :  data=30 ;
   790 :  data=30 ;
   791 :  data=35 ;
   792 :  data=13 ;
   793 :  data=-43 ;
   794 :  data=-77 ;
   795 :  data=-63 ;
   796 :  data=-77 ;
   797 :  data=-174 ;
   798 :  data=-312 ;
   799 :  data=-437 ;
   800 :  data=-493 ;
   801 :  data=-435 ;
   802 :  data=-318 ;
   803 :  data=-230 ;
   804 :  data=-156 ;
   805 :  data=-100 ;
   806 :  data=-136 ;
   807 :  data=-245 ;
   808 :  data=-361 ;
   809 :  data=-478 ;
   810 :  data=-533 ;
   811 :  data=-450 ;
   812 :  data=-338 ;
   813 :  data=-312 ;
   814 :  data=-308 ;
   815 :  data=-286 ;
   816 :  data=-329 ;
   817 :  data=-443 ;
   818 :  data=-535 ;
   819 :  data=-545 ;
   820 :  data=-501 ;
   821 :  data=-498 ;
   822 :  data=-571 ;
   823 :  data=-662 ;
   824 :  data=-794 ;
   825 :  data=-991 ;
   826 :  data=-1099 ;
   827 :  data=-1039 ;
   828 :  data=-953 ;
   829 :  data=-864 ;
   830 :  data=-692 ;
   831 :  data=-586 ;
   832 :  data=-697 ;
   833 :  data=-892 ;
   834 :  data=-1024 ;
   835 :  data=-1050 ;
   836 :  data=-912 ;
   837 :  data=-692 ;
   838 :  data=-578 ;
   839 :  data=-583 ;
   840 :  data=-647 ;
   841 :  data=-821 ;
   842 :  data=-1052 ;
   843 :  data=-1160 ;
   844 :  data=-1108 ;
   845 :  data=-1000 ;
   846 :  data=-954 ;
   847 :  data=-1038 ;
   848 :  data=-1174 ;
   849 :  data=-1250 ;
   850 :  data=-1304 ;
   851 :  data=-1347 ;
   852 :  data=-1295 ;
   853 :  data=-1213 ;
   854 :  data=-1201 ;
   855 :  data=-1166 ;
   856 :  data=-1071 ;
   857 :  data=-1017 ;
   858 :  data=-970 ;
   859 :  data=-886 ;
   860 :  data=-919 ;
   861 :  data=-1101 ;
   862 :  data=-1259 ;
   863 :  data=-1344 ;
   864 :  data=-1402 ;
   865 :  data=-1394 ;
   866 :  data=-1341 ;
   867 :  data=-1350 ;
   868 :  data=-1405 ;
   869 :  data=-1427 ;
   870 :  data=-1462 ;
   871 :  data=-1602 ;
   872 :  data=-1808 ;
   873 :  data=-1911 ;
   874 :  data=-1835 ;
   875 :  data=-1729 ;
   876 :  data=-1724 ;
   877 :  data=-1742 ;
   878 :  data=-1726 ;
   879 :  data=-1748 ;
   880 :  data=-1778 ;
   881 :  data=-1713 ;
   882 :  data=-1593 ;
   883 :  data=-1513 ;
   884 :  data=-1476 ;
   885 :  data=-1481 ;
   886 :  data=-1537 ;
   887 :  data=-1625 ;
   888 :  data=-1739 ;
   889 :  data=-1851 ;
   890 :  data=-1890 ;
   891 :  data=-1856 ;
   892 :  data=-1826 ;
   893 :  data=-1802 ;
   894 :  data=-1747 ;
   895 :  data=-1705 ;
   896 :  data=-1728 ;
   897 :  data=-1804 ;
   898 :  data=-1897 ;
   899 :  data=-1973 ;
   900 :  data=-2010 ;
   901 :  data=-2032 ;
   902 :  data=-2060 ;
   903 :  data=-2059 ;
   904 :  data=-2020 ;
   905 :  data=-2008 ;
   906 :  data=-2049 ;
   907 :  data=-2078 ;
   908 :  data=-2067 ;
   909 :  data=-2065 ;
   910 :  data=-2100 ;
   911 :  data=-2145 ;
   912 :  data=-2191 ;
   913 :  data=-2227 ;
   914 :  data=-2226 ;
   915 :  data=-2216 ;
   916 :  data=-2239 ;
   917 :  data=-2243 ;
   918 :  data=-2181 ;
   919 :  data=-2114 ;
   920 :  data=-2086 ;
   921 :  data=-2045 ;
   922 :  data=-1986 ;
   923 :  data=-1971 ;
   924 :  data=-2011 ;
   925 :  data=-2054 ;
   926 :  data=-2076 ;
   927 :  data=-2083 ;
   928 :  data=-2068 ;
   929 :  data=-2011 ;
   930 :  data=-1894 ;
   931 :  data=-1742 ;
   932 :  data=-1634 ;
   933 :  data=-1627 ;
   934 :  data=-1690 ;
   935 :  data=-1752 ;
   936 :  data=-1790 ;
   937 :  data=-1819 ;
   938 :  data=-1842 ;
   939 :  data=-1851 ;
   940 :  data=-1825 ;
   941 :  data=-1748 ;
   942 :  data=-1661 ;
   943 :  data=-1645 ;
   944 :  data=-1697 ;
   945 :  data=-1750 ;
   946 :  data=-1783 ;
   947 :  data=-1765 ;
   948 :  data=-1650 ;
   949 :  data=-1530 ;
   950 :  data=-1520 ;
   951 :  data=-1549 ;
   952 :  data=-1559 ;
   953 :  data=-1646 ;
   954 :  data=-1776 ;
   955 :  data=-1794 ;
   956 :  data=-1765 ;
   957 :  data=-1799 ;
   958 :  data=-1790 ;
   959 :  data=-1705 ;
   960 :  data=-1694 ;
   961 :  data=-1744 ;
   962 :  data=-1731 ;
   963 :  data=-1718 ;
   964 :  data=-1789 ;
   965 :  data=-1854 ;
   966 :  data=-1858 ;
   967 :  data=-1869 ;
   968 :  data=-1903 ;
   969 :  data=-1899 ;
   970 :  data=-1854 ;
   971 :  data=-1836 ;
   972 :  data=-1877 ;
   973 :  data=-1913 ;
   974 :  data=-1888 ;
   975 :  data=-1841 ;
   976 :  data=-1804 ;
   977 :  data=-1776 ;
   978 :  data=-1814 ;
   979 :  data=-1929 ;
   980 :  data=-1991 ;
   981 :  data=-1953 ;
   982 :  data=-1945 ;
   983 :  data=-1994 ;
   984 :  data=-1970 ;
   985 :  data=-1855 ;
   986 :  data=-1770 ;
   987 :  data=-1756 ;
   988 :  data=-1759 ;
   989 :  data=-1758 ;
   990 :  data=-1773 ;
   991 :  data=-1789 ;
   992 :  data=-1761 ;
   993 :  data=-1706 ;
   994 :  data=-1677 ;
   995 :  data=-1681 ;
   996 :  data=-1698 ;
   997 :  data=-1736 ;
   998 :  data=-1765 ;
   999 :  data=-1753 ;
   1000 : data=-1746 ;
   1001 : data=-1757 ;
   1002 : data=-1702 ;
   1003 : data=-1596 ;
   1004 : data=-1533 ;
   1005 : data=-1496 ;
   1006 : data=-1452 ;
   1007 : data=-1452 ;
   1008 : data=-1466 ;
   1009 : data=-1419 ;
   1010 : data=-1377 ;
   1011 : data=-1393 ;
   1012 : data=-1373 ;
   1013 : data=-1292 ;
   1014 : data=-1252 ;
   1015 : data=-1260 ;
   1016 : data=-1258 ;
   1017 : data=-1254 ;
   1018 : data=-1249 ;
   1019 : data=-1214 ;
   1020 : data=-1188 ;
   1021 : data=-1203 ;
   1022 : data=-1201 ;
   1023 : data=-1172 ;
   1024 : data=-1188 ;
   1025 : data=-1211 ;
   1026 : data=-1132 ;
   1027 : data=-1007 ;
   1028 : data=-974 ;
   1029 : data=-994 ;
   1030 : data=-955 ;
   1031 : data=-913 ;
   1032 : data=-943 ;
   1033 : data=-943 ;
   1034 : data=-834 ;
   1035 : data=-723 ;
   1036 : data=-689 ;
   1037 : data=-652 ;
   1038 : data=-565 ;
   1039 : data=-515 ;
   1040 : data=-550 ;
   1041 : data=-581 ;
   1042 : data=-524 ;
   1043 : data=-422 ;
   1044 : data=-349 ;
   1045 : data=-291 ;
   1046 : data=-202 ;
   1047 : data=-115 ;
   1048 : data=-93 ;
   1049 : data=-141 ;
   1050 : data=-227 ;
   1051 : data=-293 ;
   1052 : data=-276 ;
   1053 : data=-196 ;
   1054 : data=-152 ;
   1055 : data=-179 ;
   1056 : data=-222 ;
   1057 : data=-244 ;
   1058 : data=-234 ;
   1059 : data=-168 ;
   1060 : data=-73 ;
   1061 : data=-14 ;
   1062 : data=6 ;
   1063 : data=28 ;
   1064 : data=36 ;
   1065 : data=26 ;
   1066 : data=69 ;
   1067 : data=162 ;
   1068 : data=208 ;
   1069 : data=196 ;
   1070 : data=194 ;
   1071 : data=205 ;
   1072 : data=225 ;
   1073 : data=295 ;
   1074 : data=368 ;
   1075 : data=358 ;
   1076 : data=320 ;
   1077 : data=336 ;
   1078 : data=384 ;
   1079 : data=437 ;
   1080 : data=484 ;
   1081 : data=495 ;
   1082 : data=532 ;
   1083 : data=652 ;
   1084 : data=722 ;
   1085 : data=694 ;
   1086 : data=778 ;
   1087 : data=1003 ;
   1088 : data=1106 ;
   1089 : data=1043 ;
   1090 : data=1037 ;
   1091 : data=1136 ;
   1092 : data=1207 ;
   1093 : data=1192 ;
   1094 : data=1105 ;
   1095 : data=1010 ;
   1096 : data=1020 ;
   1097 : data=1135 ;
   1098 : data=1202 ;
   1099 : data=1145 ;
   1100 : data=1061 ;
   1101 : data=1048 ;
   1102 : data=1069 ;
   1103 : data=1033 ;
   1104 : data=959 ;
   1105 : data=949 ;
   1106 : data=1019 ;
   1107 : data=1105 ;
   1108 : data=1159 ;
   1109 : data=1135 ;
   1110 : data=1059 ;
   1111 : data=1066 ;
   1112 : data=1137 ;
   1113 : data=1081 ;
   1114 : data=950 ;
   1115 : data=981 ;
   1116 : data=1113 ;
   1117 : data=1094 ;
   1118 : data=957 ;
   1119 : data=896 ;
   1120 : data=924 ;
   1121 : data=945 ;
   1122 : data=916 ;
   1123 : data=857 ;
   1124 : data=844 ;
   1125 : data=940 ;
   1126 : data=1078 ;
   1127 : data=1134 ;
   1128 : data=1098 ;
   1129 : data=1072 ;
   1130 : data=1098 ;
   1131 : data=1102 ;
   1132 : data=1049 ;
   1133 : data=1030 ;
   1134 : data=1081 ;
   1135 : data=1098 ;
   1136 : data=1030 ;
   1137 : data=945 ;
   1138 : data=880 ;
   1139 : data=853 ;
   1140 : data=896 ;
   1141 : data=960 ;
   1142 : data=971 ;
   1143 : data=966 ;
   1144 : data=984 ;
   1145 : data=995 ;
   1146 : data=1030 ;
   1147 : data=1115 ;
   1148 : data=1154 ;
   1149 : data=1122 ;
   1150 : data=1162 ;
   1151 : data=1277 ;
   1152 : data=1296 ;
   1153 : data=1234 ;
   1154 : data=1274 ;
   1155 : data=1410 ;
   1156 : data=1503 ;
   1157 : data=1560 ;
   1158 : data=1623 ;
   1159 : data=1614 ;
   1160 : data=1544 ;
   1161 : data=1548 ;
   1162 : data=1626 ;
   1163 : data=1671 ;
   1164 : data=1710 ;
   1165 : data=1788 ;
   1166 : data=1825 ;
   1167 : data=1827 ;
   1168 : data=1864 ;
   1169 : data=1860 ;
   1170 : data=1777 ;
   1171 : data=1774 ;
   1172 : data=1881 ;
   1173 : data=1930 ;
   1174 : data=1903 ;
   1175 : data=1895 ;
   1176 : data=1854 ;
   1177 : data=1773 ;
   1178 : data=1794 ;
   1179 : data=1898 ;
   1180 : data=1906 ;
   1181 : data=1801 ;
   1182 : data=1682 ;
   1183 : data=1582 ;
   1184 : data=1541 ;
   1185 : data=1604 ;
   1186 : data=1700 ;
   1187 : data=1759 ;
   1188 : data=1825 ;
   1189 : data=1946 ;
   1190 : data=2070 ;
   1191 : data=2117 ;
   1192 : data=2064 ;
   1193 : data=1998 ;
   1194 : data=2042 ;
   1195 : data=2152 ;
   1196 : data=2180 ;
   1197 : data=2142 ;
   1198 : data=2154 ;
   1199 : data=2175 ;
               
      default:                 
            data=    'd0;     

endcase

end



endmodule





