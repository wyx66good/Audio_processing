
/*************
Author:wyx
Times :2024.7.3
hanning 1024 *256
**************/

module x_7(
        input      clk,
        input wire [9:0]i,
        output reg [8:0] data
   );

always@(posedge clk)begin
case(i)
   0 :   data= 9'd257;
   1 :   data= 9'd257;
   2 :   data= 9'd257;
   3 :   data= 9'd257;
   4 :   data= 9'd257;
   5 :   data= 9'd257;
   6 :   data= 9'd257;
   7 :   data= 9'd257;
   8 :   data= 9'd257;
   9 :   data= 9'd257;
   10 :  data= 9'd257;
   11 :  data= 9'd257;
   12 :  data= 9'd256;
   13 :  data= 9'd256;
   14 :  data= 9'd256;
   15 :  data= 9'd256;
   16 :  data= 9'd256;
   17 :  data= 9'd256;
   18 :  data= 9'd256;
   19 :  data= 9'd256;
   20 :  data= 9'd255;
   21 :  data= 9'd255;
   22 :  data= 9'd255;
   23 :  data= 9'd255;
   24 :  data= 9'd255;
   25 :  data= 9'd254;
   26 :  data= 9'd254;
   27 :  data= 9'd254;
   28 :  data= 9'd254;
   29 :  data= 9'd254;
   30 :  data= 9'd253;
   31 :  data= 9'd253;
   32 :  data= 9'd253;
   33 :  data= 9'd253;
   34 :  data= 9'd252;
   35 :  data= 9'd252;
   36 :  data= 9'd252;
   37 :  data= 9'd251;
   38 :  data= 9'd251;
   39 :  data= 9'd251;
   40 :  data= 9'd251;
   41 :  data= 9'd250;
   42 :  data= 9'd250;
   43 :  data= 9'd250;
   44 :  data= 9'd249;
   45 :  data= 9'd249;
   46 :  data= 9'd249;
   47 :  data= 9'd248;
   48 :  data= 9'd248;
   49 :  data= 9'd247;
   50 :  data= 9'd247;
   51 :  data= 9'd247;
   52 :  data= 9'd246;
   53 :  data= 9'd246;
   54 :  data= 9'd245;
   55 :  data= 9'd245;
   56 :  data= 9'd245;
   57 :  data= 9'd244;
   58 :  data= 9'd244;
   59 :  data= 9'd243;
   60 :  data= 9'd243;
   61 :  data= 9'd242;
   62 :  data= 9'd242;
   63 :  data= 9'd241;
   64 :  data= 9'd241;
   65 :  data= 9'd240;
   66 :  data= 9'd240;
   67 :  data= 9'd240;
   68 :  data= 9'd239;
   69 :  data= 9'd239;
   70 :  data= 9'd238;
   71 :  data= 9'd238;
   72 :  data= 9'd237;
   73 :  data= 9'd236;
   74 :  data= 9'd236;
   75 :  data= 9'd235;
   76 :  data= 9'd235;
   77 :  data= 9'd234;
   78 :  data= 9'd234;
   79 :  data= 9'd233;
   80 :  data= 9'd233;
   81 :  data= 9'd232;
   82 :  data= 9'd232;
   83 :  data= 9'd231;
   84 :  data= 9'd230;
   85 :  data= 9'd230;
   86 :  data= 9'd229;
   87 :  data= 9'd229;
   88 :  data= 9'd228;
   89 :  data= 9'd228;
   90 :  data= 9'd227;
   91 :  data= 9'd226;
   92 :  data= 9'd226;
   93 :  data= 9'd225;
   94 :  data= 9'd224;
   95 :  data= 9'd224;
   96 :  data= 9'd223;
   97 :  data= 9'd223;
   98 :  data= 9'd222;
   99 :  data= 9'd221;
   100 :  data=9'd221;
   101 :  data=9'd220;
   102 :  data=9'd220;
   103 :  data=9'd219;
   104 :  data=9'd218;
   105 :  data=9'd218;
   106 :  data=9'd217;
   107 :  data=9'd216;
   108 :  data=9'd216;
   109 :  data=9'd215;
   110 :  data=9'd214;
   111 :  data=9'd214;
   112 :  data=9'd213;
   113 :  data=9'd212;
   114 :  data=9'd212;
   115 :  data=9'd211;
   116 :  data=9'd210;
   117 :  data=9'd210;
   118 :  data=9'd209;
   119 :  data=9'd208;
   120 :  data=9'd208;
   121 :  data=9'd207;
   122 :  data=9'd206;
   123 :  data=9'd206;
   124 :  data=9'd205;
   125 :  data=9'd204;
   126 :  data=9'd204;
   127 :  data=9'd203;
   128 :  data=9'd202;
   129 :  data=9'd202;
   130 :  data=9'd201;
   131 :  data=9'd200;
   132 :  data=9'd200;
   133 :  data=9'd199;
   134 :  data=9'd198;
   135 :  data=9'd198;
   136 :  data=9'd197;
   137 :  data=9'd196;
   138 :  data=9'd196;
   139 :  data=9'd195;
   140 :  data=9'd194;
   141 :  data=9'd194;
   142 :  data=9'd193;
   143 :  data=9'd192;
   144 :  data=9'd192;
   145 :  data=9'd191;
   146 :  data=9'd191;
   147 :  data=9'd190;
   148 :  data=9'd189;
   149 :  data=9'd189;
   150 :  data=9'd188;
   151 :  data=9'd187;
   152 :  data=9'd187;
   153 :  data=9'd186;
   154 :  data=9'd185;
   155 :  data=9'd185;
   156 :  data=9'd184;
   157 :  data=9'd184;
   158 :  data=9'd183;
   159 :  data=9'd182;
   160 :  data=9'd182;
   161 :  data=9'd181;
   162 :  data=9'd180;
   163 :  data=9'd180;
   164 :  data=9'd179;
   165 :  data=9'd179;
   166 :  data=9'd178;
   167 :  data=9'd177;
   168 :  data=9'd177;
   169 :  data=9'd176;
   170 :  data=9'd176;
   171 :  data=9'd175;
   172 :  data=9'd175;
   173 :  data=9'd174;
   174 :  data=9'd173;
   175 :  data=9'd173;
   176 :  data=9'd172;
   177 :  data=9'd172;
   178 :  data=9'd171;
   179 :  data=9'd171;
   180 :  data=9'd170;
   181 :  data=9'd170;
   182 :  data=9'd169;
   183 :  data=9'd169;
   184 :  data=9'd168;
   185 :  data=9'd168;
   186 :  data=9'd167;
   187 :  data=9'd167;
   188 :  data=9'd166;
   189 :  data=9'd166;
   190 :  data=9'd165;
   191 :  data=9'd165;
   192 :  data=9'd164;
   193 :  data=9'd164;
   194 :  data=9'd163;
   195 :  data=9'd163;
   196 :  data=9'd162;
   197 :  data=9'd162;
   198 :  data=9'd161;
   199 :  data=9'd161;
   200 :  data=9'd161;
   201 :  data=9'd160;
   202 :  data=9'd160;
   203 :  data=9'd159;
   204 :  data=9'd159;
   205 :  data=9'd159;
   206 :  data=9'd158;
   207 :  data=9'd158;
   208 :  data=9'd157;
   209 :  data=9'd157;
   210 :  data=9'd157;
   211 :  data=9'd156;
   212 :  data=9'd156;
   213 :  data=9'd156;
   214 :  data=9'd155;
   215 :  data=9'd155;
   216 :  data=9'd155;
   217 :  data=9'd154;
   218 :  data=9'd154;
   219 :  data=9'd154;
   220 :  data=9'd153;
   221 :  data=9'd153;
   222 :  data=9'd153;
   223 :  data=9'd153;
   224 :  data=9'd152;
   225 :  data=9'd152;
   226 :  data=9'd152;
   227 :  data=9'd152;
   228 :  data=9'd151;
   229 :  data=9'd151;
   230 :  data=9'd151;
   231 :  data=9'd151;
   232 :  data=9'd151;
   233 :  data=9'd150;
   234 :  data=9'd150;
   235 :  data=9'd150;
   236 :  data=9'd150;
   237 :  data=9'd150;
   238 :  data=9'd150;
   239 :  data=9'd150;
   240 :  data=9'd149;
   241 :  data=9'd149;
   242 :  data=9'd149;
   243 :  data=9'd149;
   244 :  data=9'd149;
   245 :  data=9'd149;
   246 :  data=9'd149;
   247 :  data=9'd149;
   248 :  data=9'd149;
   249 :  data=9'd149;
   250 :  data=9'd149;
   251 :  data=9'd148;
   252 :  data=9'd148;
   253 :  data=9'd148;
   254 :  data=9'd148;
   255 :  data=9'd148;
   256 :  data=9'd148;
   257 :  data=9'd148;
   258 :  data=9'd148;
   259 :  data=9'd148;
   260 :  data=9'd148;
   261 :  data=9'd149;
   262 :  data=9'd149;
   263 :  data=9'd149;
   264 :  data=9'd149;
   265 :  data=9'd149;
   266 :  data=9'd149;
   267 :  data=9'd149;
   268 :  data=9'd149;
   269 :  data=9'd149;
   270 :  data=9'd149;
   271 :  data=9'd149;
   272 :  data=9'd150;
   273 :  data=9'd150;
   274 :  data=9'd150;
   275 :  data=9'd150;
   276 :  data=9'd150;
   277 :  data=9'd150;
   278 :  data=9'd150;
   279 :  data=9'd151;
   280 :  data=9'd151;
   281 :  data=9'd151;
   282 :  data=9'd151;
   283 :  data=9'd151;
   284 :  data=9'd152;
   285 :  data=9'd152;
   286 :  data=9'd152;
   287 :  data=9'd152;
   288 :  data=9'd153;
   289 :  data=9'd153;
   290 :  data=9'd153;
   291 :  data=9'd153;
   292 :  data=9'd154;
   293 :  data=9'd154;
   294 :  data=9'd154;
   295 :  data=9'd155;
   296 :  data=9'd155;
   297 :  data=9'd155;
   298 :  data=9'd156;
   299 :  data=9'd156;
   300 :  data=9'd156;
   301 :  data=9'd157;
   302 :  data=9'd157;
   303 :  data=9'd157;
   304 :  data=9'd158;
   305 :  data=9'd158;
   306 :  data=9'd159;
   307 :  data=9'd159;
   308 :  data=9'd159;
   309 :  data=9'd160;
   310 :  data=9'd160;
   311 :  data=9'd161;
   312 :  data=9'd161;
   313 :  data=9'd161;
   314 :  data=9'd162;
   315 :  data=9'd162;
   316 :  data=9'd163;
   317 :  data=9'd163;
   318 :  data=9'd164;
   319 :  data=9'd164;
   320 :  data=9'd165;
   321 :  data=9'd165;
   322 :  data=9'd166;
   323 :  data=9'd166;
   324 :  data=9'd167;
   325 :  data=9'd167;
   326 :  data=9'd168;
   327 :  data=9'd168;
   328 :  data=9'd169;
   329 :  data=9'd169;
   330 :  data=9'd170;
   331 :  data=9'd170;
   332 :  data=9'd171;
   333 :  data=9'd171;
   334 :  data=9'd172;
   335 :  data=9'd172;
   336 :  data=9'd173;
   337 :  data=9'd173;
   338 :  data=9'd174;
   339 :  data=9'd175;
   340 :  data=9'd175;
   341 :  data=9'd176;
   342 :  data=9'd176;
   343 :  data=9'd177;
   344 :  data=9'd177;
   345 :  data=9'd178;
   346 :  data=9'd179;
   347 :  data=9'd179;
   348 :  data=9'd180;
   349 :  data=9'd180;
   350 :  data=9'd181;
   351 :  data=9'd182;
   352 :  data=9'd182;
   353 :  data=9'd183;
   354 :  data=9'd184;
   355 :  data=9'd184;
   356 :  data=9'd185;
   357 :  data=9'd185;
   358 :  data=9'd186;
   359 :  data=9'd187;
   360 :  data=9'd187;
   361 :  data=9'd188;
   362 :  data=9'd189;
   363 :  data=9'd189;
   364 :  data=9'd190;
   365 :  data=9'd191;
   366 :  data=9'd191;
   367 :  data=9'd192;
   368 :  data=9'd192;
   369 :  data=9'd193;
   370 :  data=9'd194;
   371 :  data=9'd194;
   372 :  data=9'd195;
   373 :  data=9'd196;
   374 :  data=9'd196;
   375 :  data=9'd197;
   376 :  data=9'd198;
   377 :  data=9'd198;
   378 :  data=9'd199;
   379 :  data=9'd200;
   380 :  data=9'd200;
   381 :  data=9'd201;
   382 :  data=9'd202;
   383 :  data=9'd202;
   384 :  data=9'd203;
   385 :  data=9'd204;
   386 :  data=9'd204;
   387 :  data=9'd205;
   388 :  data=9'd206;
   389 :  data=9'd206;
   390 :  data=9'd207;
   391 :  data=9'd208;
   392 :  data=9'd208;
   393 :  data=9'd209;
   394 :  data=9'd210;
   395 :  data=9'd210;
   396 :  data=9'd211;
   397 :  data=9'd212;
   398 :  data=9'd212;
   399 :  data=9'd213;
   400 :  data=9'd214;
   401 :  data=9'd214;
   402 :  data=9'd215;
   403 :  data=9'd216;
   404 :  data=9'd216;
   405 :  data=9'd217;
   406 :  data=9'd218;
   407 :  data=9'd218;
   408 :  data=9'd219;
   409 :  data=9'd220;
   410 :  data=9'd220;
   411 :  data=9'd221;
   412 :  data=9'd221;
   413 :  data=9'd222;
   414 :  data=9'd223;
   415 :  data=9'd223;
   416 :  data=9'd224;
   417 :  data=9'd224;
   418 :  data=9'd225;
   419 :  data=9'd226;
   420 :  data=9'd226;
   421 :  data=9'd227;
   422 :  data=9'd228;
   423 :  data=9'd228;
   424 :  data=9'd229;
   425 :  data=9'd229;
   426 :  data=9'd230;
   427 :  data=9'd230;
   428 :  data=9'd231;
   429 :  data=9'd232;
   430 :  data=9'd232;
   431 :  data=9'd233;
   432 :  data=9'd233;
   433 :  data=9'd234;
   434 :  data=9'd234;
   435 :  data=9'd235;
   436 :  data=9'd235;
   437 :  data=9'd236;
   438 :  data=9'd236;
   439 :  data=9'd237;
   440 :  data=9'd238;
   441 :  data=9'd238;
   442 :  data=9'd239;
   443 :  data=9'd239;
   444 :  data=9'd240;
   445 :  data=9'd240;
   446 :  data=9'd240;
   447 :  data=9'd241;
   448 :  data=9'd241;
   449 :  data=9'd242;
   450 :  data=9'd242;
   451 :  data=9'd243;
   452 :  data=9'd243;
   453 :  data=9'd244;
   454 :  data=9'd244;
   455 :  data=9'd245;
   456 :  data=9'd245;
   457 :  data=9'd245;
   458 :  data=9'd246;
   459 :  data=9'd246;
   460 :  data=9'd247;
   461 :  data=9'd247;
   462 :  data=9'd247;
   463 :  data=9'd248;
   464 :  data=9'd248;
   465 :  data=9'd249;
   466 :  data=9'd249;
   467 :  data=9'd249;
   468 :  data=9'd250;
   469 :  data=9'd250;
   470 :  data=9'd250;
   471 :  data=9'd251;
   472 :  data=9'd251;
   473 :  data=9'd251;
   474 :  data=9'd251;
   475 :  data=9'd252;
   476 :  data=9'd252;
   477 :  data=9'd252;
   478 :  data=9'd253;
   479 :  data=9'd253;
   480 :  data=9'd253;
   481 :  data=9'd253;
   482 :  data=9'd254;
   483 :  data=9'd254;
   484 :  data=9'd254;
   485 :  data=9'd254;
   486 :  data=9'd254;
   487 :  data=9'd255;
   488 :  data=9'd255;
   489 :  data=9'd255;
   490 :  data=9'd255;
   491 :  data=9'd255;
   492 :  data=9'd256;
   493 :  data=9'd256;
   494 :  data=9'd256;
   495 :  data=9'd256;
   496 :  data=9'd256;
   497 :  data=9'd256;
   498 :  data=9'd256;
   499 :  data=9'd256;
   500 :  data=9'd257;
   501 :  data=9'd257;
   502 :  data=9'd257;
   503 :  data=9'd257;
   504 :  data=9'd257;
   505 :  data=9'd257;
   506 :  data=9'd257;
   507 :  data=9'd257;
   508 :  data=9'd257;
   509 :  data=9'd257;
   510 :  data=9'd257;
   511 :  data=9'd257;
   512 :  data=9'd257;
   513 :  data=9'd257;
   514 :  data=9'd257;
   515 :  data=9'd257;
   516 :  data=9'd257;
   517 :  data=9'd257;
   518 :  data=9'd257;
   519 :  data=9'd257;
   520 :  data=9'd257;
   521 :  data=9'd257;
   522 :  data=9'd257;
   523 :  data=9'd257;
   524 :  data=9'd256;
   525 :  data=9'd256;
   526 :  data=9'd256;
   527 :  data=9'd256;
   528 :  data=9'd256;
   529 :  data=9'd256;
   530 :  data=9'd256;
   531 :  data=9'd256;
   532 :  data=9'd255;
   533 :  data=9'd255;
   534 :  data=9'd255;
   535 :  data=9'd255;
   536 :  data=9'd255;
   537 :  data=9'd254;
   538 :  data=9'd254;
   539 :  data=9'd254;
   540 :  data=9'd254;
   541 :  data=9'd254;
   542 :  data=9'd253;
   543 :  data=9'd253;
   544 :  data=9'd253;
   545 :  data=9'd253;
   546 :  data=9'd252;
   547 :  data=9'd252;
   548 :  data=9'd252;
   549 :  data=9'd251;
   550 :  data=9'd251;
   551 :  data=9'd251;
   552 :  data=9'd251;
   553 :  data=9'd250;
   554 :  data=9'd250;
   555 :  data=9'd250;
   556 :  data=9'd249;
   557 :  data=9'd249;
   558 :  data=9'd249;
   559 :  data=9'd248;
   560 :  data=9'd248;
   561 :  data=9'd247;
   562 :  data=9'd247;
   563 :  data=9'd247;
   564 :  data=9'd246;
   565 :  data=9'd246;
   566 :  data=9'd245;
   567 :  data=9'd245;
   568 :  data=9'd245;
   569 :  data=9'd244;
   570 :  data=9'd244;
   571 :  data=9'd243;
   572 :  data=9'd243;
   573 :  data=9'd242;
   574 :  data=9'd242;
   575 :  data=9'd241;
   576 :  data=9'd241;
   577 :  data=9'd240;
   578 :  data=9'd240;
   579 :  data=9'd240;
   580 :  data=9'd239;
   581 :  data=9'd239;
   582 :  data=9'd238;
   583 :  data=9'd238;
   584 :  data=9'd237;
   585 :  data=9'd236;
   586 :  data=9'd236;
   587 :  data=9'd235;
   588 :  data=9'd235;
   589 :  data=9'd234;
   590 :  data=9'd234;
   591 :  data=9'd233;
   592 :  data=9'd233;
   593 :  data=9'd232;
   594 :  data=9'd232;
   595 :  data=9'd231;
   596 :  data=9'd230;
   597 :  data=9'd230;
   598 :  data=9'd229;
   599 :  data=9'd229;
   600 :  data=9'd228;
   601 :  data=9'd228;
   602 :  data=9'd227;
   603 :  data=9'd226;
   604 :  data=9'd226;
   605 :  data=9'd225;
   606 :  data=9'd224;
   607 :  data=9'd224;
   608 :  data=9'd223;
   609 :  data=9'd223;
   610 :  data=9'd222;
   611 :  data=9'd221;
   612 :  data=9'd221;
   613 :  data=9'd220;
   614 :  data=9'd220;
   615 :  data=9'd219;
   616 :  data=9'd218;
   617 :  data=9'd218;
   618 :  data=9'd217;
   619 :  data=9'd216;
   620 :  data=9'd216;
   621 :  data=9'd215;
   622 :  data=9'd214;
   623 :  data=9'd214;
   624 :  data=9'd213;
   625 :  data=9'd212;
   626 :  data=9'd212;
   627 :  data=9'd211;
   628 :  data=9'd210;
   629 :  data=9'd210;
   630 :  data=9'd209;
   631 :  data=9'd208;
   632 :  data=9'd208;
   633 :  data=9'd207;
   634 :  data=9'd206;
   635 :  data=9'd206;
   636 :  data=9'd205;
   637 :  data=9'd204;
   638 :  data=9'd204;
   639 :  data=9'd203;
   640 :  data=9'd202;
   641 :  data=9'd202;
   642 :  data=9'd201;
   643 :  data=9'd200;
   644 :  data=9'd200;
   645 :  data=9'd199;
   646 :  data=9'd198;
   647 :  data=9'd198;
   648 :  data=9'd197;
   649 :  data=9'd196;
   650 :  data=9'd196;
   651 :  data=9'd195;
   652 :  data=9'd194;
   653 :  data=9'd194;
   654 :  data=9'd193;
   655 :  data=9'd192;
   656 :  data=9'd192;
   657 :  data=9'd191;
   658 :  data=9'd191;
   659 :  data=9'd190;
   660 :  data=9'd189;
   661 :  data=9'd189;
   662 :  data=9'd188;
   663 :  data=9'd187;
   664 :  data=9'd187;
   665 :  data=9'd186;
   666 :  data=9'd185;
   667 :  data=9'd185;
   668 :  data=9'd184;
   669 :  data=9'd184;
   670 :  data=9'd183;
   671 :  data=9'd182;
   672 :  data=9'd182;
   673 :  data=9'd181;
   674 :  data=9'd180;
   675 :  data=9'd180;
   676 :  data=9'd179;
   677 :  data=9'd179;
   678 :  data=9'd178;
   679 :  data=9'd177;
   680 :  data=9'd177;
   681 :  data=9'd176;
   682 :  data=9'd176;
   683 :  data=9'd175;
   684 :  data=9'd175;
   685 :  data=9'd174;
   686 :  data=9'd173;
   687 :  data=9'd173;
   688 :  data=9'd172;
   689 :  data=9'd172;
   690 :  data=9'd171;
   691 :  data=9'd171;
   692 :  data=9'd170;
   693 :  data=9'd170;
   694 :  data=9'd169;
   695 :  data=9'd169;
   696 :  data=9'd168;
   697 :  data=9'd168;
   698 :  data=9'd167;
   699 :  data=9'd167;
   700 :  data=9'd166;
   701 :  data=9'd166;
   702 :  data=9'd165;
   703 :  data=9'd165;
   704 :  data=9'd164;
   705 :  data=9'd164;
   706 :  data=9'd163;
   707 :  data=9'd163;
   708 :  data=9'd162;
   709 :  data=9'd162;
   710 :  data=9'd161;
   711 :  data=9'd161;
   712 :  data=9'd161;
   713 :  data=9'd160;
   714 :  data=9'd160;
   715 :  data=9'd159;
   716 :  data=9'd159;
   717 :  data=9'd159;
   718 :  data=9'd158;
   719 :  data=9'd158;
   720 :  data=9'd157;
   721 :  data=9'd157;
   722 :  data=9'd157;
   723 :  data=9'd156;
   724 :  data=9'd156;
   725 :  data=9'd156;
   726 :  data=9'd155;
   727 :  data=9'd155;
   728 :  data=9'd155;
   729 :  data=9'd154;
   730 :  data=9'd154;
   731 :  data=9'd154;
   732 :  data=9'd153;
   733 :  data=9'd153;
   734 :  data=9'd153;
   735 :  data=9'd153;
   736 :  data=9'd152;
   737 :  data=9'd152;
   738 :  data=9'd152;
   739 :  data=9'd152;
   740 :  data=9'd151;
   741 :  data=9'd151;
   742 :  data=9'd151;
   743 :  data=9'd151;
   744 :  data=9'd151;
   745 :  data=9'd150;
   746 :  data=9'd150;
   747 :  data=9'd150;
   748 :  data=9'd150;
   749 :  data=9'd150;
   750 :  data=9'd150;
   751 :  data=9'd150;
   752 :  data=9'd149;
   753 :  data=9'd149;
   754 :  data=9'd149;
   755 :  data=9'd149;
   756 :  data=9'd149;
   757 :  data=9'd149;
   758 :  data=9'd149;
   759 :  data=9'd149;
   760 :  data=9'd149;
   761 :  data=9'd149;
   762 :  data=9'd149;
   763 :  data=9'd148;
   764 :  data=9'd148;
   765 :  data=9'd148;
   766 :  data=9'd148;
   767 :  data=9'd148;
   768 :  data=9'd148;
   769 :  data=9'd148;
   770 :  data=9'd148;
   771 :  data=9'd148;
   772 :  data=9'd148;
   773 :  data=9'd149;
   774 :  data=9'd149;
   775 :  data=9'd149;
   776 :  data=9'd149;
   777 :  data=9'd149;
   778 :  data=9'd149;
   779 :  data=9'd149;
   780 :  data=9'd149;
   781 :  data=9'd149;
   782 :  data=9'd149;
   783 :  data=9'd149;
   784 :  data=9'd150;
   785 :  data=9'd150;
   786 :  data=9'd150;
   787 :  data=9'd150;
   788 :  data=9'd150;
   789 :  data=9'd150;
   790 :  data=9'd150;
   791 :  data=9'd151;
   792 :  data=9'd151;
   793 :  data=9'd151;
   794 :  data=9'd151;
   795 :  data=9'd151;
   796 :  data=9'd152;
   797 :  data=9'd152;
   798 :  data=9'd152;
   799 :  data=9'd152;
   800 :  data=9'd153;
   801 :  data=9'd153;
   802 :  data=9'd153;
   803 :  data=9'd153;
   804 :  data=9'd154;
   805 :  data=9'd154;
   806 :  data=9'd154;
   807 :  data=9'd155;
   808 :  data=9'd155;
   809 :  data=9'd155;
   810 :  data=9'd156;
   811 :  data=9'd156;
   812 :  data=9'd156;
   813 :  data=9'd157;
   814 :  data=9'd157;
   815 :  data=9'd157;
   816 :  data=9'd158;
   817 :  data=9'd158;
   818 :  data=9'd159;
   819 :  data=9'd159;
   820 :  data=9'd159;
   821 :  data=9'd160;
   822 :  data=9'd160;
   823 :  data=9'd161;
   824 :  data=9'd161;
   825 :  data=9'd161;
   826 :  data=9'd162;
   827 :  data=9'd162;
   828 :  data=9'd163;
   829 :  data=9'd163;
   830 :  data=9'd164;
   831 :  data=9'd164;
   832 :  data=9'd165;
   833 :  data=9'd165;
   834 :  data=9'd166;
   835 :  data=9'd166;
   836 :  data=9'd167;
   837 :  data=9'd167;
   838 :  data=9'd168;
   839 :  data=9'd168;
   840 :  data=9'd169;
   841 :  data=9'd169;
   842 :  data=9'd170;
   843 :  data=9'd170;
   844 :  data=9'd171;
   845 :  data=9'd171;
   846 :  data=9'd172;
   847 :  data=9'd172;
   848 :  data=9'd173;
   849 :  data=9'd173;
   850 :  data=9'd174;
   851 :  data=9'd175;
   852 :  data=9'd175;
   853 :  data=9'd176;
   854 :  data=9'd176;
   855 :  data=9'd177;
   856 :  data=9'd177;
   857 :  data=9'd178;
   858 :  data=9'd179;
   859 :  data=9'd179;
   860 :  data=9'd180;
   861 :  data=9'd180;
   862 :  data=9'd181;
   863 :  data=9'd182;
   864 :  data=9'd182;
   865 :  data=9'd183;
   866 :  data=9'd184;
   867 :  data=9'd184;
   868 :  data=9'd185;
   869 :  data=9'd185;
   870 :  data=9'd186;
   871 :  data=9'd187;
   872 :  data=9'd187;
   873 :  data=9'd188;
   874 :  data=9'd189;
   875 :  data=9'd189;
   876 :  data=9'd190;
   877 :  data=9'd191;
   878 :  data=9'd191;
   879 :  data=9'd192;
   880 :  data=9'd192;
   881 :  data=9'd193;
   882 :  data=9'd194;
   883 :  data=9'd194;
   884 :  data=9'd195;
   885 :  data=9'd196;
   886 :  data=9'd196;
   887 :  data=9'd197;
   888 :  data=9'd198;
   889 :  data=9'd198;
   890 :  data=9'd199;
   891 :  data=9'd200;
   892 :  data=9'd200;
   893 :  data=9'd201;
   894 :  data=9'd202;
   895 :  data=9'd202;
   896 :  data=9'd203;
   897 :  data=9'd204;
   898 :  data=9'd204;
   899 :  data=9'd205;
   900 :  data=9'd206;
   901 :  data=9'd206;
   902 :  data=9'd207;
   903 :  data=9'd208;
   904 :  data=9'd208;
   905 :  data=9'd209;
   906 :  data=9'd210;
   907 :  data=9'd210;
   908 :  data=9'd211;
   909 :  data=9'd212;
   910 :  data=9'd212;
   911 :  data=9'd213;
   912 :  data=9'd214;
   913 :  data=9'd214;
   914 :  data=9'd215;
   915 :  data=9'd216;
   916 :  data=9'd216;
   917 :  data=9'd217;
   918 :  data=9'd218;
   919 :  data=9'd218;
   920 :  data=9'd219;
   921 :  data=9'd220;
   922 :  data=9'd220;
   923 :  data=9'd221;
   924 :  data=9'd221;
   925 :  data=9'd222;
   926 :  data=9'd223;
   927 :  data=9'd223;
   928 :  data=9'd224;
   929 :  data=9'd224;
   930 :  data=9'd225;
   931 :  data=9'd226;
   932 :  data=9'd226;
   933 :  data=9'd227;
   934 :  data=9'd228;
   935 :  data=9'd228;
   936 :  data=9'd229;
   937 :  data=9'd229;
   938 :  data=9'd230;
   939 :  data=9'd230;
   940 :  data=9'd231;
   941 :  data=9'd232;
   942 :  data=9'd232;
   943 :  data=9'd233;
   944 :  data=9'd233;
   945 :  data=9'd234;
   946 :  data=9'd234;
   947 :  data=9'd235;
   948 :  data=9'd235;
   949 :  data=9'd236;
   950 :  data=9'd236;
   951 :  data=9'd237;
   952 :  data=9'd238;
   953 :  data=9'd238;
   954 :  data=9'd239;
   955 :  data=9'd239;
   956 :  data=9'd240;
   957 :  data=9'd240;
   958 :  data=9'd240;
   959 :  data=9'd241;
   960 :  data=9'd241;
   961 :  data=9'd242;
   962 :  data=9'd242;
   963 :  data=9'd243;
   964 :  data=9'd243;
   965 :  data=9'd244;
   966 :  data=9'd244;
   967 :  data=9'd245;
   968 :  data=9'd245;
   969 :  data=9'd245;
   970 :  data=9'd246;
   971 :  data=9'd246;
   972 :  data=9'd247;
   973 :  data=9'd247;
   974 :  data=9'd247;
   975 :  data=9'd248;
   976 :  data=9'd248;
   977 :  data=9'd249;
   978 :  data=9'd249;
   979 :  data=9'd249;
   980 :  data=9'd250;
   981 :  data=9'd250;
   982 :  data=9'd250;
   983 :  data=9'd251;
   984 :  data=9'd251;
   985 :  data=9'd251;
   986 :  data=9'd251;
   987 :  data=9'd252;
   988 :  data=9'd252;
   989 :  data=9'd252;
   990 :  data=9'd253;
   991 :  data=9'd253;
   992 :  data=9'd253;
   993 :  data=9'd253;
   994 :  data=9'd254;
   995 :  data=9'd254;
   996 :  data=9'd254;
   997 :  data=9'd254;
   998 :  data=9'd254;
   999 :  data=9'd255;
   1000 : data=9'd255;
   1001 : data=9'd255;
   1002 : data=9'd255;
   1003 : data=9'd255;
   1004 : data=9'd256;
   1005 : data=9'd256;
   1006 : data=9'd256;
   1007 : data=9'd256;
   1008 : data=9'd256;
   1009 : data=9'd256;
   1010 : data=9'd256;
   1011 : data=9'd256;
   1012 : data=9'd257;
   1013 : data=9'd257;
   1014 : data=9'd257;
   1015 : data=9'd257;
   1016 : data=9'd257;
   1017 : data=9'd257;
   1018 : data=9'd257;
   1019 : data=9'd257;
   1020 : data=9'd257;
   1021 : data=9'd257;
   1022 : data=9'd257;
   1023 : data=9'd257;
                  
      default:                 
            data=    'd0;     

endcase

end






endmodule