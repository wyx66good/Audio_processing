/*************
Author:wyx
Times :2024.5.30
���ҷ��ȵ��� ������128
**************/


module sin_Amplitude_modulation(
        input wire [9:0]i,
        output reg [7:0] data
   );


always @(*) begin
case(i)
   0 :   data= 0    ;
   1 :   data= 1    ;
   2 :   data= 2    ;
   3 :   data= 4    ;
   4 :   data= 5    ;
   5 :   data= 6    ;
   6 :   data= 8    ;
   7 :   data= 9    ;
   8 :   data= 10   ;
   9 :   data= 12   ;
   10 :  data= 13   ;
   11 :  data= 14   ;
   12 :  data= 16   ;
   13 :  data= 17   ;
   14 :  data= 18   ;
   15 :  data= 20   ;
   16 :  data= 21   ;
   17 :  data= 22   ;
   18 :  data= 23   ;
   19 :  data= 25   ;
   20 :  data= 26   ;
   21 :  data= 27   ;
   22 :  data= 29   ;
   23 :  data= 30   ;
   24 :  data= 31   ;
   25 :  data= 33   ;
   26 :  data= 34   ;
   27 :  data= 35   ;
   28 :  data= 36   ;
   29 :  data= 38   ;
   30 :  data= 39   ;
   31 :  data= 40   ;
   32 :  data= 42   ;
   33 :  data= 43   ;
   34 :  data= 44   ;
   35 :  data= 45   ;
   36 :  data= 47   ;
   37 :  data= 48   ;
   38 :  data= 49   ;
   39 :  data= 50   ;
   40 :  data= 52   ;
   41 :  data= 53   ;
   42 :  data= 54   ;
   43 :  data= 55   ;
   44 :  data= 56   ;
   45 :  data= 58   ;
   46 :  data= 59   ;
   47 :  data= 60   ;
   48 :  data= 61   ;
   49 :  data= 62   ;
   50 :  data= 64   ;
   51 :  data= 65   ;
   52 :  data= 66   ;
   53 :  data= 67   ;
   54 :  data= 68   ;
   55 :  data= 69   ;
   56 :  data= 70   ;
   57 :  data= 71   ;
   58 :  data= 73   ;
   59 :  data= 74   ;
   60 :  data= 75   ;
   61 :  data= 76   ;
   62 :  data= 77   ;
   63 :  data= 78   ;
   64 :  data= 79   ;
   65 :  data= 80   ;
   66 :  data= 81   ;
   67 :  data= 82   ;
   68 :  data= 83   ;
   69 :  data= 84   ;
   70 :  data= 85   ;
   71 :  data= 86   ;
   72 :  data= 87   ;
   73 :  data= 88   ;
   74 :  data= 89   ;
   75 :  data= 90   ;
   76 :  data= 91   ;
   77 :  data= 92   ;
   78 :  data= 93   ;
   79 :  data= 94   ;
   80 :  data= 95   ;
   81 :  data= 96   ;
   82 :  data= 96   ;
   83 :  data= 97   ;
   84 :  data= 98   ;
   85 :  data= 99   ;
   86 :  data= 100  ;
   87 :  data= 101  ;
   88 :  data= 101  ;
   89 :  data= 102  ;
   90 :  data= 103  ;
   91 :  data= 104  ;
   92 :  data= 105  ;
   93 :  data= 105  ;
   94 :  data= 106  ;
   95 :  data= 107  ;
   96 :  data= 108  ;
   97 :  data= 108  ;
   98 :  data= 109  ;
   99 :  data= 110  ;
   100 :  data=110  ;
   101 :  data=111  ;
   102 :  data=112  ;
   103 :  data=112  ;
   104 :  data=113  ;
   105 :  data=114  ;
   106 :  data=114  ;
   107 :  data=115  ;
   108 :  data=115  ;
   109 :  data=116  ;
   110 :  data=116  ;
   111 :  data=117  ;
   112 :  data=117  ;
   113 :  data=118  ;
   114 :  data=119  ;
   115 :  data=119  ;
   116 :  data=119  ;
   117 :  data=120  ;
   118 :  data=120  ;
   119 :  data=121  ;
   120 :  data=121  ;
   121 :  data=122  ;
   122 :  data=122  ;
   123 :  data=122  ;
   124 :  data=123  ;
   125 :  data=123  ;
   126 :  data=123  ;
   127 :  data=124  ;
   128 :  data=124  ;
   129 :  data=124  ;
   130 :  data=125  ;
   131 :  data=125  ;
   132 :  data=125  ;
   133 :  data=125  ;
   134 :  data=126  ;
   135 :  data=126  ;
   136 :  data=126  ;
   137 :  data=126  ;
   138 :  data=126  ;
   139 :  data=127  ;
   140 :  data=127  ;
   141 :  data=127  ;
   142 :  data=127  ;
   143 :  data=127  ;
   144 :  data=127  ;
   145 :  data=127  ;
   146 :  data=127  ;
   147 :  data=127  ;
   148 :  data=127  ;
   149 :  data=127  ;
   150 :  data=128  ;
   151 :  data=127  ;
   152 :  data=127  ;
   153 :  data=127  ;
   154 :  data=127  ;
   155 :  data=127  ;
   156 :  data=127  ;
   157 :  data=127  ;
   158 :  data=127  ;
   159 :  data=127  ;
   160 :  data=127  ;
   161 :  data=127  ;
   162 :  data=126  ;
   163 :  data=126  ;
   164 :  data=126  ;
   165 :  data=126  ;
   166 :  data=126  ;
   167 :  data=125  ;
   168 :  data=125  ;
   169 :  data=125  ;
   170 :  data=125  ;
   171 :  data=124  ;
   172 :  data=124  ;
   173 :  data=124  ;
   174 :  data=123  ;
   175 :  data=123  ;
   176 :  data=123  ;
   177 :  data=122  ;
   178 :  data=122  ;
   179 :  data=122  ;
   180 :  data=121  ;
   181 :  data=122  ;
   182 :  data=122  ;
   183 :  data=122  ;
   184 :  data=123  ;
   185 :  data=123  ;
   186 :  data=123  ;
   187 :  data=124  ;
   188 :  data=124  ;
   189 :  data=124  ;
   190 :  data=125  ;
   191 :  data=125  ;
   192 :  data=125  ;
   193 :  data=125  ;
   194 :  data=126  ;
   195 :  data=126  ;
   196 :  data=126  ;
   197 :  data=126  ;
   198 :  data=126  ;
   199 :  data=127  ;
   200 :  data=127  ;
   201 :  data=127  ;
   202 :  data=127  ;
   203 :  data=127  ;
   204 :  data=127  ;
   205 :  data=127  ;
   206 :  data=127  ;
   207 :  data=127  ;
   208 :  data=127  ;
   209 :  data=127  ;
   210 :  data=128  ;
   211 :  data=127  ;
   212 :  data=127  ;
   213 :  data=127  ;
   214 :  data=127  ;
   215 :  data=127  ;
   216 :  data=127  ;
   217 :  data=127  ;
   218 :  data=127  ;
   219 :  data=127  ;
   220 :  data=127  ;
   221 :  data=127  ;
   222 :  data=126  ;
   223 :  data=126  ;
   224 :  data=126  ;
   225 :  data=126  ;
   226 :  data=126  ;
   227 :  data=125  ;
   228 :  data=125  ;
   229 :  data=125  ;
   230 :  data=125  ;
   231 :  data=124  ;
   232 :  data=124  ;
   233 :  data=124  ;
   234 :  data=123  ;
   235 :  data=123  ;
   236 :  data=123  ;
   237 :  data=122  ;
   238 :  data=122  ;
   239 :  data=122  ;
   240 :  data=121  ;
   241 :  data=122  ;
   242 :  data=122  ;
   243 :  data=122  ;
   244 :  data=123  ;
   245 :  data=123  ;
   246 :  data=123  ;
   247 :  data=124  ;
   248 :  data=124  ;
   249 :  data=124  ;
   250 :  data=125  ;
   251 :  data=125  ;
   252 :  data=125  ;
   253 :  data=125  ;
   254 :  data=126  ;
   255 :  data=126  ;
   256 :  data=126  ;
   257 :  data=126  ;
   258 :  data=126  ;
   259 :  data=127  ;
   260 :  data=127  ;
   261 :  data=127  ;
   262 :  data=127  ;
   263 :  data=127  ;
   264 :  data=127  ;
   265 :  data=127  ;
   266 :  data=127  ;
   267 :  data=127  ;
   268 :  data=127  ;
   269 :  data=127  ;
   270 :  data=128  ;
   271 :  data=127  ;
   272 :  data=127  ;
   273 :  data=127  ;
   274 :  data=127  ;
   275 :  data=127  ;
   276 :  data=127  ;
   277 :  data=127  ;
   278 :  data=127  ;
   279 :  data=127  ;
   280 :  data=127  ;
   281 :  data=127  ;
   282 :  data=126  ;
   283 :  data=126  ;
   284 :  data=126  ;
   285 :  data=126  ;
   286 :  data=126  ;
   287 :  data=125  ;
   288 :  data=125  ;
   289 :  data=125  ;
   290 :  data=125  ;
   291 :  data=124  ;
   292 :  data=124  ;
   293 :  data=124  ;
   294 :  data=123  ;
   295 :  data=123  ;
   296 :  data=123  ;
   297 :  data=122  ;
   298 :  data=122  ;
   299 :  data=122  ;
  300 :  data= 121  ;
   301 :  data=122  ;
   302 :  data=122  ;
   303 :  data=122  ;
   304 :  data=123  ;
   305 :  data=123  ;
   306 :  data=123  ;
   307 :  data=124  ;
   308 :  data=124  ;
   309 :  data=124  ;
   310 :  data=125  ;
   311 :  data=125  ;
   312 :  data=125  ;
   313 :  data=125  ;
   314 :  data=126  ;
   315 :  data=126  ;
   316 :  data=126  ;
   317 :  data=126  ;
   318 :  data=126  ;
   319 :  data=127  ;
   320 :  data=127  ;
   321 :  data=127  ;
   322 :  data=127  ;
   323 :  data=127  ;
   324 :  data=127  ;
   325 :  data=127  ;
   326 :  data=127  ;
   327 :  data=127  ;
   328 :  data=127  ;
   329 :  data=127  ;
   330 :  data=128  ;
   331 :  data=127  ;
   332 :  data=127  ;
   333 :  data=127  ;
   334 :  data=127  ;
   335 :  data=127  ;
   336 :  data=127  ;
   337 :  data=127  ;
   338 :  data=127  ;
   339 :  data=127  ;
   340 :  data=127  ;
   341 :  data=127  ;
   342 :  data=126  ;
   343 :  data=126  ;
   344 :  data=126  ;
   345 :  data=126  ;
   346 :  data=126  ;
   347 :  data=125  ;
   348 :  data=125  ;
   349 :  data=125  ;
   350 :  data=125  ;
   351 :  data=124  ;
   352 :  data=124  ;
   353 :  data=124  ;
   354 :  data=123  ;
   355 :  data=123  ;
   356 :  data=123  ;
   357 :  data=122  ;
   358 :  data=122  ;
   359 :  data=122  ;
   360 :  data=121  ;
   361 :  data=122  ;
   362 :  data=122  ;
   363 :  data=122  ;
   364 :  data=123  ;
   365 :  data=123  ;
   366 :  data=123  ;
   367 :  data=124  ;
   368 :  data=124  ;
   369 :  data=124  ;
   370 :  data=125  ;
   371 :  data=125  ;
   372 :  data=125  ;
   373 :  data=125  ;
   374 :  data=126  ;
   375 :  data=126  ;
   376 :  data=126  ;
   377 :  data=126  ;
   378 :  data=126  ;
   379 :  data=127  ;
   380 :  data=127  ;
   381 :  data=127  ;
   382 :  data=127  ;
   383 :  data=127  ;
   384 :  data=127  ;
   385 :  data=127  ;
   386 :  data=127  ;
   387 :  data=127  ;
   388 :  data=127  ;
   389 :  data=127  ;
   390 :  data=128  ;
   391 :  data=127  ;
   392 :  data=127  ;
   393 :  data=127  ;
   394 :  data=127  ;
   395 :  data=127  ;
   396 :  data=127  ;
   397 :  data=127  ;
   398 :  data=127  ;
   399 :  data=127  ;
   400 :  data=127  ;
   401 :  data=127  ;
   402 :  data=126  ;
   403 :  data=126  ;
   404 :  data=126  ;
   405 :  data=126  ;
   406 :  data=126  ;
   407 :  data=125  ;
   408 :  data=125  ;
   409 :  data=125  ;
   410 :  data=125  ;
   411 :  data=124  ;
   412 :  data=124  ;
   413 :  data=124  ;
   414 :  data=123  ;
   415 :  data=123  ;
   416 :  data=123  ;
   417 :  data=122  ;
   418 :  data=122  ;
   419 :  data=122  ;
   420 :  data=121  ;
   421 :  data=122  ;
   422 :  data=122  ;
   423 :  data=122  ;
   424 :  data=123  ;
   425 :  data=123  ;
   426 :  data=123  ;
   427 :  data=124  ;
   428 :  data=124  ;
   429 :  data=124  ;
   430 :  data=125  ;
   431 :  data=125  ;
   432 :  data=125  ;
   433 :  data=125  ;
   434 :  data=126  ;
   435 :  data=126  ;
   436 :  data=126  ;
   437 :  data=126  ;
   438 :  data=126  ;
   439 :  data=127  ;
   440 :  data=127  ;
   441 :  data=127  ;
   442 :  data=127  ;
   443 :  data=127  ;
   444 :  data=127  ;
   445 :  data=127  ;
   446 :  data=127  ;
   447 :  data=127  ;
   448 :  data=127  ;
   449 :  data=127  ;
   450 :  data=128  ;
   451 :  data=127  ;
   452 :  data=127  ;
   453 :  data=127  ;
   454 :  data=127  ;
   455 :  data=127  ;
   456 :  data=127  ;
   457 :  data=127  ;
   458 :  data=127  ;
   459 :  data=127  ;
   460 :  data=127  ;
   461 :  data=127  ;
   462 :  data=126  ;
   463 :  data=126  ;
   464 :  data=126  ;
   465 :  data=126  ;
   466 :  data=126  ;
   467 :  data=125  ;
   468 :  data=125  ;
   469 :  data=125  ;
   470 :  data=125  ;
   471 :  data=124  ;
   472 :  data=124  ;
   473 :  data=124  ;
   474 :  data=123  ;
   475 :  data=123  ;
   476 :  data=123  ;
   477 :  data=122  ;
   478 :  data=122  ;
   479 :  data=122  ;
   480 :  data=121  ;
   481 :  data=121  ;
   482 :  data=120  ;
   483 :  data=120  ;
   484 :  data=119  ;
   485 :  data=119  ;
   486 :  data=119  ;
   487 :  data=118  ;
   488 :  data=117  ;
   489 :  data=117  ;
   490 :  data=116  ;
   491 :  data=116  ;
   492 :  data=115  ;
   493 :  data=115  ;
   494 :  data=114  ;
   495 :  data=114  ;
   496 :  data=113  ;
   497 :  data=112  ;
   498 :  data=112  ;
   499 :  data=111  ;
   500 :  data=110  ;
   501 :  data=110  ;
   502 :  data=109  ;
   503 :  data=108  ;
   504 :  data=108  ;
   505 :  data=107  ;
   506 :  data=106  ;
   507 :  data=105  ;
   508 :  data=105  ;
   509 :  data=104  ;
   510 :  data=103  ;
   511 :  data=102  ;
   512 :  data=101  ;
   513 :  data=101  ;
   514 :  data=100  ;
   515 :  data=99   ;
   516 :  data=98   ;
   517 :  data=97   ;
   518 :  data=96   ;
   519 :  data=96   ;
   520 :  data=95   ;
   521 :  data=94   ;
   522 :  data=93   ;
   523 :  data=92   ;
   524 :  data=91   ;
   525 :  data=90   ;
   526 :  data=89   ;
   527 :  data=88   ;
   528 :  data=87   ;
   529 :  data=86   ;
   530 :  data=85   ;
   531 :  data=84   ;
   532 :  data=83   ;
   533 :  data=82   ;
   534 :  data=81   ;
   535 :  data=80   ;
   536 :  data=79   ;
   537 :  data=78   ;
   538 :  data=77   ;
   539 :  data=76   ;
   540 :  data=75   ;
   541 :  data=74   ;
   542 :  data=73   ;
   543 :  data=71   ;
   544 :  data=70   ;
   545 :  data=69   ;
   546 :  data=68   ;
   547 :  data=67   ;
   548 :  data=66   ;
   549 :  data=65   ;
   550 :  data=64   ;
   551 :  data=62   ;
   552 :  data=61   ;
   553 :  data=60   ;
   554 :  data=59   ;
   555 :  data=58   ;
   556 :  data=56   ;
   557 :  data=55   ;
   558 :  data=54   ;
   559 :  data=53   ;
   560 :  data=52   ;
   561 :  data=50   ;
   562 :  data=49   ;
   563 :  data=48   ;
   564 :  data=47   ;
   565 :  data=45   ;
   566 :  data=44   ;
   567 :  data=43   ;
   568 :  data=42   ;
   569 :  data=40   ;
   570 :  data=39   ;
   571 :  data=38   ;
   572 :  data=36   ;
   573 :  data=35   ;
   574 :  data=34   ;
   575 :  data=33   ;
   576 :  data=31   ;
   577 :  data=30   ;
   578 :  data=29   ;
   579 :  data=27   ;
   580 :  data=26   ;
   581 :  data=25   ;
   582 :  data=23   ;
   583 :  data=22   ;
   584 :  data=21   ;
   585 :  data=20   ;
   586 :  data=18   ;
   587 :  data=17   ;
   588 :  data=16   ;
   589 :  data=14   ;
   590 :  data=13   ;
   591 :  data=12   ;
   592 :  data=10   ;
   593 :  data=9    ;
   594 :  data=8    ;
   595 :  data=6    ;
   596 :  data=5    ;
   597 :  data=4    ;
   598 :  data=2    ;
   599 :  data=1    ;
               
      default:                 
            data=    'd0;     

endcase

end



endmodule



