`timescale 1ns/1ns
module hpss_fir
#(
    parameter DATA_WIDTH = 16,
    parameter FILTER_ORDER = 100
)
(
    input                       sck,
    input                       rst_n,

    output reg [DATA_WIDTH - 1:0]  ldata,
    output reg [DATA_WIDTH - 1:0]  rdata,

    input   [DATA_WIDTH - 1:0]  data,
    input                       r_vld,
    input                       l_vld
);

parameter signed [15:0] b [0:FILTER_ORDER] = {
   16'sd72,   // 0.00221 * 2^15
    16'sd56,   // 0.00170 * 2^15
    16'sd25,   // 0.00076 * 2^15
    -16'sd16,   // -0.00048 * 2^15
    -16'sd58,   // -0.00178 * 2^15
    -16'sd94,   // -0.00288 * 2^15
    -16'sd112,   // -0.00343 * 2^15
    -16'sd104,   // -0.00317 * 2^15
    -16'sd64,   // -0.00195 * 2^15
    16'sd4,   // 0.00013 * 2^15
    16'sd88,   // 0.00269 * 2^15
    16'sd168,   // 0.00512 * 2^15
    16'sd219,   // 0.00667 * 2^15
    16'sd219,   // 0.00669 * 2^15
    16'sd158,   // 0.00482 * 2^15
    16'sd39,   // 0.00118 * 2^15
    -16'sd117,   // -0.00356 * 2^15
    -16'sd270,   // -0.00825 * 2^15
    -16'sd379,   // -0.01156 * 2^15
    -16'sd403,   // -0.01230 * 2^15
    -16'sd321,   // -0.00981 * 2^15
    -16'sd139,   // -0.00424 * 2^15
    16'sd109,   // 0.00333 * 2^15
    16'sd365,   // 0.01114 * 2^15
    16'sd560,   // 0.01708 * 2^15
    16'sd632,   // 0.01928 * 2^15
    16'sd546,   // 0.01667 * 2^15
    16'sd307,   // 0.00937 * 2^15
    -16'sd39,   // -0.00120 * 2^15
    -16'sd412,   // -0.01258 * 2^15
    -16'sd716,   // -0.02184 * 2^15
    -16'sd863,   // -0.02633 * 2^15
    -16'sd801,   // -0.02445 * 2^15
    -16'sd529,   // -0.01615 * 2^15
    -16'sd101,   // -0.00309 * 2^15
    16'sd383,   // 0.01170 * 2^15
    16'sd803,   // 0.02451 * 2^15
    16'sd1046,   // 0.03192 * 2^15
    16'sd1039,   // 0.03170 * 2^15
    16'sd770,   // 0.02351 * 2^15
    16'sd296,   // 0.00904 * 2^15
    -16'sd272,   // -0.00831 * 2^15
    -16'sd795,   // -0.02425 * 2^15
    -16'sd1137,   // -0.03470 * 2^15
    -16'sd1208,   // -0.03685 * 2^15
    -16'sd981,   // -0.02994 * 2^15
    -16'sd508,   // -0.01549 * 2^15
    16'sd99,   // 0.00301 * 2^15
    16'sd688,   // 0.02100 * 2^15
    16'sd1114,   // 0.03399 * 2^15
    16'sd1269,   // 0.03871 * 2^15
    16'sd1114,   // 0.03399 * 2^15
    16'sd688,   // 0.02100 * 2^15
    16'sd99,   // 0.00301 * 2^15
    -16'sd508,   // -0.01549 * 2^15
    -16'sd981,   // -0.02994 * 2^15
    -16'sd1208,   // -0.03685 * 2^15
    -16'sd1137,   // -0.03470 * 2^15
    -16'sd795,   // -0.02425 * 2^15
    -16'sd272,   // -0.00831 * 2^15
    16'sd296,   // 0.00904 * 2^15
    16'sd770,   // 0.02351 * 2^15
    16'sd1039,   // 0.03170 * 2^15
    16'sd1046,   // 0.03192 * 2^15
    16'sd803,   // 0.02451 * 2^15
    16'sd383,   // 0.01170 * 2^15
    -16'sd101,   // -0.00309 * 2^15
    -16'sd529,   // -0.01615 * 2^15
    -16'sd801,   // -0.02445 * 2^15
    -16'sd863,   // -0.02633 * 2^15
    -16'sd716,   // -0.02184 * 2^15
    -16'sd412,   // -0.01258 * 2^15
    -16'sd39,   // -0.00120 * 2^15
    16'sd307,   // 0.00937 * 2^15
    16'sd546,   // 0.01667 * 2^15
    16'sd632,   // 0.01928 * 2^15
    16'sd560,   // 0.01708 * 2^15
    16'sd365,   // 0.01114 * 2^15
    16'sd109,   // 0.00333 * 2^15
    -16'sd139,   // -0.00424 * 2^15
    -16'sd321,   // -0.00981 * 2^15
    -16'sd403,   // -0.01230 * 2^15
    -16'sd379,   // -0.01156 * 2^15
    -16'sd270,   // -0.00825 * 2^15
    -16'sd117,   // -0.00356 * 2^15
    16'sd39,   // 0.00118 * 2^15
    16'sd158,   // 0.00482 * 2^15
    16'sd219,   // 0.00669 * 2^15
    16'sd219,   // 0.00667 * 2^15
    16'sd168,   // 0.00512 * 2^15
    16'sd88,   // 0.00269 * 2^15
    16'sd4,   // 0.00013 * 2^15
    -16'sd64,   // -0.00195 * 2^15
    -16'sd104,   // -0.00317 * 2^15
    -16'sd112,   // -0.00343 * 2^15
    -16'sd94,   // -0.00288 * 2^15
    -16'sd58,   // -0.00178 * 2^15
    -16'sd16,   // -0.00048 * 2^15
    16'sd25,   // 0.00076 * 2^15
    16'sd56,   // 0.00170 * 2^15
    16'sd72   // 0.00221 * 2^15
};


reg signed [DATA_WIDTH - 1:0] x_left [0:FILTER_ORDER];  
reg signed [DATA_WIDTH - 1:0] x_right [0:FILTER_ORDER]; 


reg signed [31:0] acc_left;
reg signed [31:0] acc_right;

integer i;

reg  [5:0]                 cnt_2000k;
    always @(posedge sck or negedge rst_n)
    begin
    	if(~rst_n)
    	    cnt_2000k <= 6'h0;
    	else
    	begin
    		if(cnt_2000k == 6'd6)
    		    cnt_2000k <= 6'h0;
    		else
    		    cnt_2000k <= cnt_2000k + 1'b1;
    	end
    end


//always @(posedge sck or negedge rst_n)
//begin
//    if(~rst_n)
//    begin
//        ldata <= {DATA_WIDTH{1'b0}};
//        for (i = 0; i <= FILTER_ORDER; i = i + 1)
//            x_left[i] <= {DATA_WIDTH{1'b0}};
//    end
//    else if(l_vld && cnt_2000k == 6'd6)
//    begin
//
//        for (i = FILTER_ORDER; i > 0; i = i - 1)
//            x_left[i] <= x_left[i - 1];
//        x_left[0] <= data;
//
//
//        acc_left = 0;
//        for (i = 0; i <= FILTER_ORDER; i = i + 1)
//            acc_left = acc_left + x_left[i] * b[i];
//
//        ldata <= acc_left[31:16]*3; 
//end
//     else
//         ldata <=  ldata;
//    
//end


always @(posedge sck or negedge rst_n)
begin
    if(~rst_n)
    begin
        rdata <= {DATA_WIDTH{1'b0}};
        for (i = 0; i <= FILTER_ORDER; i = i + 1)
            x_right[i] <= {DATA_WIDTH{1'b0}};
    end
    else if(r_vld && cnt_2000k == 6'd6)
    begin

        for (i = FILTER_ORDER; i > 0; i = i - 1)
            x_right[i] <= x_right[i - 1];
        x_right[0] <= data;


        acc_right = 0;
        for (i = 0; i <= FILTER_ORDER; i = i + 1)
            acc_right = acc_right + x_right[i] * b[i];

        rdata <= acc_right[31:16]*3; 
end
     else
      rdata  <=  rdata;
    
end

endmodule // i2s_loop
