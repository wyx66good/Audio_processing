
/*************
Author:wyx
Times :2024.7.3
hanning_1024 *256
**************/

module hanning(
        input      clk,
        input wire [9:0]i,
        output reg [7:0] data
   );

always@(posedge clk)begin
case(i)
   0 :   data= 8'd0    ;
   1 :   data= 8'd0    ;
   2 :   data= 8'd0    ;
   3 :   data= 8'd0    ;
   4 :   data= 8'd10    ;
   5 :   data= 8'd10    ;
   6 :   data= 8'd10    ;
   7 :   data= 8'd10    ;
   8 :   data= 8'd10    ;
   9 :   data= 8'd10    ;
   10 :  data= 8'd20    ;
   11 :  data= 8'd20    ;
   12 :  data= 8'd20    ;
   13 :  data= 8'd20    ;
   14 :  data= 8'd20    ;
   15 :  data= 8'd20    ;
   16 :  data= 8'd21    ;
   17 :  data= 8'd21    ;
   18 :  data= 8'd21    ;
   19 :  data= 8'd21    ;
   20 :  data= 8'd21    ;
   21 :  data= 8'd21    ;
   22 :  data= 8'd21    ;
   23 :  data= 8'd21    ;
   24 :  data= 8'd21    ;
   25 :  data= 8'd21    ;
   26 :  data= 8'd21    ;
   27 :  data= 8'd22    ;
   28 :  data= 8'd22    ;
   29 :  data= 8'd22    ;
   30 :  data= 8'd22    ;
   31 :  data= 8'd22    ;
   32 :  data= 8'd22    ;
   33 :  data= 8'd22    ;
   34 :  data= 8'd23    ;
   35 :  data= 8'd23    ;
   36 :  data= 8'd23    ;
   37 :  data= 8'd23    ;
   38 :  data= 8'd23    ;
   39 :  data= 8'd23    ;
   40 :  data= 8'd24    ;
   41 :  data= 8'd24    ;
   42 :  data= 8'd24    ;
   43 :  data= 8'd24    ;
   44 :  data= 8'd24    ;
   45 :  data= 8'd24    ;
   46 :  data= 8'd25    ;
   47 :  data= 8'd25    ;
   48 :  data= 8'd25    ;
   49 :  data= 8'd25    ;
   50 :  data= 8'd25    ;
   51 :  data= 8'd26    ;
   52 :  data= 8'd26    ;
   53 :  data= 8'd26    ;
   54 :  data= 8'd26    ;
   55 :  data= 8'd27    ;
   56 :  data= 8'd27    ;
   57 :  data= 8'd27    ;
   58 :  data= 8'd27    ;
   59 :  data= 8'd28    ;
   60 :  data= 8'd28    ;
   61 :  data= 8'd28    ;
   62 :  data= 8'd28    ;
   63 :  data= 8'd29    ;
   64 :  data= 8'd29    ;
   65 :  data= 8'd29    ;
   66 :  data= 8'd30    ;
   67 :  data= 8'd30    ;
   68 :  data= 8'd30    ;
   69 :  data= 8'd30    ;
   70 :  data= 8'd31    ;
   71 :  data= 8'd31    ;
   72 :  data= 8'd31    ;
   73 :  data= 8'd32    ;
   74 :  data= 8'd32    ;
   75 :  data= 8'd32    ;
   76 :  data= 8'd33    ;
   77 :  data= 8'd33    ;
   78 :  data= 8'd33    ;
   79 :  data= 8'd34    ;
   80 :  data= 8'd34    ;
   81 :  data= 8'd34    ;
   82 :  data= 8'd35    ;
   83 :  data= 8'd35    ;
   84 :  data= 8'd35    ;
   85 :  data= 8'd36    ;
   86 :  data= 8'd36    ;
   87 :  data= 8'd36    ;
   88 :  data= 8'd37    ;
   89 :  data= 8'd37    ;
   90 :  data= 8'd38    ;
   91 :  data= 8'd38    ;
   92 :  data= 8'd38    ;
   93 :  data= 8'd39    ;
   94 :  data= 8'd39    ;
   95 :  data= 8'd39    ;
   96 :  data= 8'd40    ;
   97 :  data= 8'd40    ;
   98 :  data= 8'd41    ;
   99 :  data= 8'd41    ;
   100 :  data=8'd42    ;
   101 :  data=8'd42    ;
   102 :  data=8'd42    ;
   103 :  data=8'd43    ;
   104 :  data=8'd43    ;
   105 :  data=8'd44    ;
   106 :  data=8'd44    ;
   107 :  data=8'd45    ;
   108 :  data=8'd45    ;
   109 :  data=8'd45    ;
   110 :  data=8'd46    ;
   111 :  data=8'd46    ;
   112 :  data=8'd47    ;
   113 :  data=8'd47    ;
   114 :  data=8'd48    ;
   115 :  data=8'd48    ;
   116 :  data=8'd49    ;
   117 :  data=8'd49    ;
   118 :  data=8'd50    ;
   119 :  data=8'd50    ;
   120 :  data=8'd51    ;
   121 :  data=8'd51    ;
   122 :  data=8'd52    ;
   123 :  data=8'd52    ;
   124 :  data=8'd53    ;
   125 :  data=8'd53    ;
   126 :  data=8'd54    ;
   127 :  data=8'd54    ;
   128 :  data=8'd55    ;
   129 :  data=8'd55    ;
   130 :  data=8'd56    ;
   131 :  data=8'd56    ;
   132 :  data=8'd57    ;
   133 :  data=8'd57    ;
   134 :  data=8'd58    ;
   135 :  data=8'd58    ;
   136 :  data=8'd59    ;
   137 :  data=8'd59    ;
   138 :  data=8'd60    ;
   139 :  data=8'd60    ;
   140 :  data=8'd61    ;
   141 :  data=8'd61    ;
   142 :  data=8'd62    ;
   143 :  data=8'd63    ;
   144 :  data=8'd63    ;
   145 :  data=8'd64    ;
   146 :  data=8'd64    ;
   147 :  data=8'd65    ;
   148 :  data=8'd65    ;
   149 :  data=8'd66    ;
   150 :  data=8'd67    ;
   151 :  data=8'd67    ;
   152 :  data=8'd68    ;
   153 :  data=8'd68    ;
   154 :  data=8'd69    ;
   155 :  data=8'd69    ;
   156 :  data=8'd70    ;
   157 :  data=8'd71    ;
   158 :  data=8'd71    ;
   159 :  data=8'd72    ;
   160 :  data=8'd72    ;
   161 :  data=8'd73    ;
   162 :  data=8'd74    ;
   163 :  data=8'd74    ;
   164 :  data=8'd75    ;
   165 :  data=8'd75    ;
   166 :  data=8'd76    ;
   167 :  data=8'd77    ;
   168 :  data=8'd77    ;
   169 :  data=8'd78    ;
   170 :  data=8'd79    ;
   171 :  data=8'd79    ;
   172 :  data=8'd80    ;
   173 :  data=8'd80    ;
   174 :  data=8'd81    ;
   175 :  data=8'd82    ;
   176 :  data=8'd82    ;
   177 :  data=8'd83    ;
   178 :  data=8'd84    ;
   179 :  data=8'd84    ;
   180 :  data=8'd85    ;
   181 :  data=8'd86    ;
   182 :  data=8'd86    ;
   183 :  data=8'd87    ;
   184 :  data=8'd88    ;
   185 :  data=8'd88    ;
   186 :  data=8'd89    ;
   187 :  data=8'd89    ;
   188 :  data=8'd90    ;
   189 :  data=8'd91    ;
   190 :  data=8'd91    ;
   191 :  data=8'd92    ;
   192 :  data=8'd93    ;
   193 :  data=8'd93    ;
   194 :  data=8'd94    ;
   195 :  data=8'd95    ;
   196 :  data=8'd95    ;
   197 :  data=8'd96    ;
   198 :  data=8'd97    ;
   199 :  data=8'd98    ;
   200 :  data=8'd98    ;
   201 :  data=8'd99    ;
   202 :  data=8'd100   ;
   203 :  data=8'd100   ;
   204 :  data=8'd101   ;
   205 :  data=8'd102   ;
   206 :  data=8'd102   ;
   207 :  data=8'd103   ;
   208 :  data=8'd104   ;
   209 :  data=8'd104   ;
   210 :  data=8'd105   ;
   211 :  data=8'd106   ;
   212 :  data=8'd106   ;
   213 :  data=8'd107   ;
   214 :  data=8'd108   ;
   215 :  data=8'd109   ;
   216 :  data=8'd109   ;
   217 :  data=8'd110   ;
   218 :  data=8'd111   ;
   219 :  data=8'd111   ;
   220 :  data=8'd112   ;
   221 :  data=8'd113   ;
   222 :  data=8'd114   ;
   223 :  data=8'd114   ;
   224 :  data=8'd115   ;
   225 :  data=8'd116   ;
   226 :  data=8'd116   ;
   227 :  data=8'd117   ;
   228 :  data=8'd118   ;
   229 :  data=8'd118   ;
   230 :  data=8'd119   ;
   231 :  data=8'd120   ;
   232 :  data=8'd121   ;
   233 :  data=8'd121   ;
   234 :  data=8'd122   ;
   235 :  data=8'd123   ;
   236 :  data=8'd123   ;
   237 :  data=8'd124   ;
   238 :  data=8'd125   ;
   239 :  data=8'd126   ;
   240 :  data=8'd126   ;
   241 :  data=8'd127   ;
   242 :  data=8'd128   ;
   243 :  data=8'd129   ;
   244 :  data=8'd129   ;
   245 :  data=8'd130   ;
   246 :  data=8'd131   ;
   247 :  data=8'd131   ;
   248 :  data=8'd132   ;
   249 :  data=8'd133   ;
   250 :  data=8'd134   ;
   251 :  data=8'd134   ;
   252 :  data=8'd135   ;
   253 :  data=8'd136   ;
   254 :  data=8'd136   ;
   255 :  data=8'd137   ;
   256 :  data=8'd138   ;
   257 :  data=8'd139   ;
   258 :  data=8'd139   ;
   259 :  data=8'd140   ;
   260 :  data=8'd141   ;
   261 :  data=8'd142   ;
   262 :  data=8'd142   ;
   263 :  data=8'd143   ;
   264 :  data=8'd144   ;
   265 :  data=8'd144   ;
   266 :  data=8'd145   ;
   267 :  data=8'd146   ;
   268 :  data=8'd147   ;
   269 :  data=8'd147   ;
   270 :  data=8'd148   ;
   271 :  data=8'd149   ;
   272 :  data=8'd149   ;
   273 :  data=8'd150   ;
   274 :  data=8'd151   ;
   275 :  data=8'd152   ;
   276 :  data=8'd152   ;
   277 :  data=8'd153   ;
   278 :  data=8'd154   ;
   279 :  data=8'd154   ;
   280 :  data=8'd155   ;
   281 :  data=8'd156   ;
   282 :  data=8'd157   ;
   283 :  data=8'd157   ;
   284 :  data=8'd158   ;
   285 :  data=8'd159   ;
   286 :  data=8'd159   ;
   287 :  data=8'd160   ;
   288 :  data=8'd161   ;
   289 :  data=8'd162   ;
   290 :  data=8'd162   ;
   291 :  data=8'd163   ;
   292 :  data=8'd164   ;
   293 :  data=8'd164   ;
   294 :  data=8'd165   ;
   295 :  data=8'd166   ;
   296 :  data=8'd167   ;
   297 :  data=8'd167   ;
   298 :  data=8'd168   ;
   299 :  data=8'd169   ;
   300 :  data=8'd169   ;
   301 :  data=8'd170   ;
   302 :  data=8'd171   ;
   303 :  data=8'd171   ;
   304 :  data=8'd172   ;
   305 :  data=8'd173   ;
   306 :  data=8'd174   ;
   307 :  data=8'd174   ;
   308 :  data=8'd175   ;
   309 :  data=8'd176   ;
   310 :  data=8'd176   ;
   311 :  data=8'd177   ;
   312 :  data=8'd178   ;
   313 :  data=8'd178   ;
   314 :  data=8'd179   ;
   315 :  data=8'd180   ;
   316 :  data=8'd180   ;
   317 :  data=8'd181   ;
   318 :  data=8'd182   ;
   319 :  data=8'd182   ;
   320 :  data=8'd183   ;
   321 :  data=8'd184   ;
   322 :  data=8'd184   ;
   323 :  data=8'd185   ;
   324 :  data=8'd186   ;
   325 :  data=8'd186   ;
   326 :  data=8'd187   ;
   327 :  data=8'd188   ;
   328 :  data=8'd188   ;
   329 :  data=8'd189   ;
   330 :  data=8'd190   ;
   331 :  data=8'd190   ;
   332 :  data=8'd191   ;
   333 :  data=8'd192   ;
   334 :  data=8'd192   ;
   335 :  data=8'd193   ;
   336 :  data=8'd193   ;
   337 :  data=8'd194   ;
   338 :  data=8'd195   ;
   339 :  data=8'd195   ;
   340 :  data=8'd196   ;
   341 :  data=8'd197   ;
   342 :  data=8'd197   ;
   343 :  data=8'd198   ;
   344 :  data=8'd198   ;
   345 :  data=8'd199   ;
   346 :  data=8'd200   ;
   347 :  data=8'd200   ;
   348 :  data=8'd201   ;
   349 :  data=8'd202   ;
   350 :  data=8'd202   ;
   351 :  data=8'd203   ;
   352 :  data=8'd203   ;
   353 :  data=8'd204   ;
   354 :  data=8'd205   ;
   355 :  data=8'd205   ;
   356 :  data=8'd206   ;
   357 :  data=8'd206   ;
   358 :  data=8'd207   ;
   359 :  data=8'd208   ;
   360 :  data=8'd208   ;
   361 :  data=8'd209   ;
   362 :  data=8'd209   ;
   363 :  data=8'd210   ;
   364 :  data=8'd210   ;
   365 :  data=8'd211   ;
   366 :  data=8'd212   ;
   367 :  data=8'd212   ;
   368 :  data=8'd213   ;
   369 :  data=8'd213   ;
   370 :  data=8'd214   ;
   371 :  data=8'd214   ;
   372 :  data=8'd215   ;
   373 :  data=8'd215   ;
   374 :  data=8'd216   ;
   375 :  data=8'd216   ;
   376 :  data=8'd217   ;
   377 :  data=8'd218   ;
   378 :  data=8'd218   ;
   379 :  data=8'd219   ;
   380 :  data=8'd219   ;
   381 :  data=8'd220   ;
   382 :  data=8'd220   ;
   383 :  data=8'd221   ;
   384 :  data=8'd221   ;
   385 :  data=8'd222   ;
   386 :  data=8'd222   ;
   387 :  data=8'd223   ;
   388 :  data=8'd223   ;
   389 :  data=8'd224   ;
   390 :  data=8'd224   ;
   391 :  data=8'd225   ;
   392 :  data=8'd225   ;
   393 :  data=8'd226   ;
   394 :  data=8'd226   ;
   395 :  data=8'd227   ;
   396 :  data=8'd227   ;
   397 :  data=8'd228   ;
   398 :  data=8'd228   ;
   399 :  data=8'd228   ;
   400 :  data=8'd229   ;
   401 :  data=8'd229   ;
   402 :  data=8'd230   ;
   403 :  data=8'd230   ;
   404 :  data=8'd231   ;
   405 :  data=8'd231   ;
   406 :  data=8'd232   ;
   407 :  data=8'd232   ;
   408 :  data=8'd232   ;
   409 :  data=8'd233   ;
   410 :  data=8'd233   ;
   411 :  data=8'd234   ;
   412 :  data=8'd234   ;
   413 :  data=8'd235   ;
   414 :  data=8'd235   ;
   415 :  data=8'd235   ;
   416 :  data=8'd236   ;
   417 :  data=8'd236   ;
   418 :  data=8'd237   ;
   419 :  data=8'd237   ;
   420 :  data=8'd237   ;
   421 :  data=8'd238   ;
   422 :  data=8'd238   ;
   423 :  data=8'd239   ;
   424 :  data=8'd239   ;
   425 :  data=8'd239   ;
   426 :  data=8'd240   ;
   427 :  data=8'd240   ;
   428 :  data=8'd240   ;
   429 :  data=8'd241   ;
   430 :  data=8'd241   ;
   431 :  data=8'd241   ;
   432 :  data=8'd242   ;
   433 :  data=8'd242   ;
   434 :  data=8'd242   ;
   435 :  data=8'd243   ;
   436 :  data=8'd243   ;
   437 :  data=8'd243   ;
   438 :  data=8'd244   ;
   439 :  data=8'd244   ;
   440 :  data=8'd244   ;
   441 :  data=8'd245   ;
   442 :  data=8'd245   ;
   443 :  data=8'd245   ;
   444 :  data=8'd246   ;
   445 :  data=8'd246   ;
   446 :  data=8'd246   ;
   447 :  data=8'd246   ;
   448 :  data=8'd247   ;
   449 :  data=8'd247   ;
   450 :  data=8'd247   ;
   451 :  data=8'd247   ;
   452 :  data=8'd248   ;
   453 :  data=8'd248   ;
   454 :  data=8'd248   ;
   455 :  data=8'd248   ;
   456 :  data=8'd249   ;
   457 :  data=8'd249   ;
   458 :  data=8'd249   ;
   459 :  data=8'd249   ;
   460 :  data=8'd250   ;
   461 :  data=8'd250   ;
   462 :  data=8'd250   ;
   463 :  data=8'd250   ;
   464 :  data=8'd251   ;
   465 :  data=8'd251   ;
   466 :  data=8'd251   ;
   467 :  data=8'd251   ;
   468 :  data=8'd251   ;
   469 :  data=8'd252   ;
   470 :  data=8'd252   ;
   471 :  data=8'd252   ;
   472 :  data=8'd252   ;
   473 :  data=8'd252   ;
   474 :  data=8'd252   ;
   475 :  data=8'd253   ;
   476 :  data=8'd253   ;
   477 :  data=8'd253   ;
   478 :  data=8'd253   ;
   479 :  data=8'd253   ;
   480 :  data=8'd253   ;
   481 :  data=8'd253   ;
   482 :  data=8'd254   ;
   483 :  data=8'd254   ;
   484 :  data=8'd254   ;
   485 :  data=8'd254   ;
   486 :  data=8'd254   ;
   487 :  data=8'd254   ;
   488 :  data=8'd254   ;
   489 :  data=8'd254   ;
   490 :  data=8'd254   ;
   491 :  data=8'd255   ;
   492 :  data=8'd255   ;
   493 :  data=8'd255   ;
   494 :  data=8'd255   ;
   495 :  data=8'd255   ;
   496 :  data=8'd255   ;
   497 :  data=8'd255   ;
   498 :  data=8'd255   ;
   499 :  data=8'd255   ;
   500 :  data=8'd255   ;
   501 :  data=8'd255   ;
   502 :  data=8'd255   ;
   503 :  data=8'd255   ;
   504 :  data=8'd255   ;
   505 :  data=8'd255   ;
   506 :  data=8'd255   ;
   507 :  data=8'd255   ;
   508 :  data=8'd255   ;
   509 :  data=8'd255   ;
   510 :  data=8'd255   ;
   511 :  data=8'd255   ;
   512 :  data=8'd255   ;
   513 :  data=8'd255   ;
   514 :  data=8'd255   ;
   515 :  data=8'd255   ;
   516 :  data=8'd255   ;
   517 :  data=8'd255   ;
   518 :  data=8'd255   ;
   519 :  data=8'd255   ;
   520 :  data=8'd255   ;
   521 :  data=8'd255   ;
   522 :  data=8'd255   ;
   523 :  data=8'd255   ;
   524 :  data=8'd255   ;
   525 :  data=8'd255   ;
   526 :  data=8'd255   ;
   527 :  data=8'd255   ;
   528 :  data=8'd255   ;
   529 :  data=8'd255   ;
   530 :  data=8'd255   ;
   531 :  data=8'd255   ;
   532 :  data=8'd255   ;
   533 :  data=8'd254   ;
   534 :  data=8'd254   ;
   535 :  data=8'd254   ;
   536 :  data=8'd254   ;
   537 :  data=8'd254   ;
   538 :  data=8'd254   ;
   539 :  data=8'd254   ;
   540 :  data=8'd254   ;
   541 :  data=8'd254   ;
   542 :  data=8'd253   ;
   543 :  data=8'd253   ;
   544 :  data=8'd253   ;
   545 :  data=8'd253   ;
   546 :  data=8'd253   ;
   547 :  data=8'd253   ;
   548 :  data=8'd253   ;
   549 :  data=8'd252   ;
   550 :  data=8'd252   ;
   551 :  data=8'd252   ;
   552 :  data=8'd252   ;
   553 :  data=8'd252   ;
   554 :  data=8'd252   ;
   555 :  data=8'd251   ;
   556 :  data=8'd251   ;
   557 :  data=8'd251   ;
   558 :  data=8'd251   ;
   559 :  data=8'd251   ;
   560 :  data=8'd250   ;
   561 :  data=8'd250   ;
   562 :  data=8'd250   ;
   563 :  data=8'd250   ;
   564 :  data=8'd249   ;
   565 :  data=8'd249   ;
   566 :  data=8'd249   ;
   567 :  data=8'd249   ;
   568 :  data=8'd248   ;
   569 :  data=8'd248   ;
   570 :  data=8'd248   ;
   571 :  data=8'd248   ;
   572 :  data=8'd247   ;
   573 :  data=8'd247   ;
   574 :  data=8'd247   ;
   575 :  data=8'd247   ;
   576 :  data=8'd246   ;
   577 :  data=8'd246   ;
   578 :  data=8'd246   ;
   579 :  data=8'd246   ;
   580 :  data=8'd245   ;
   581 :  data=8'd245   ;
   582 :  data=8'd245   ;
   583 :  data=8'd244   ;
   584 :  data=8'd244   ;
   585 :  data=8'd244   ;
   586 :  data=8'd243   ;
   587 :  data=8'd243   ;
   588 :  data=8'd243   ;
   589 :  data=8'd242   ;
   590 :  data=8'd242   ;
   591 :  data=8'd242   ;
   592 :  data=8'd241   ;
   593 :  data=8'd241   ;
   594 :  data=8'd241   ;
   595 :  data=8'd240   ;
   596 :  data=8'd240   ;
   597 :  data=8'd240   ;
   598 :  data=8'd239   ;
   599 :  data=8'd239   ;
   600 :  data=8'd239   ;
   601 :  data=8'd238   ;
   602 :  data=8'd238   ;
   603 :  data=8'd237   ;
   604 :  data=8'd237   ;
   605 :  data=8'd237   ;
   606 :  data=8'd236   ;
   607 :  data=8'd236   ;
   608 :  data=8'd235   ;
   609 :  data=8'd235   ;
   610 :  data=8'd235   ;
   611 :  data=8'd234   ;
   612 :  data=8'd234   ;
   613 :  data=8'd233   ;
   614 :  data=8'd233   ;
   615 :  data=8'd232   ;
   616 :  data=8'd232   ;
   617 :  data=8'd232   ;
   618 :  data=8'd231   ;
   619 :  data=8'd231   ;
   620 :  data=8'd230   ;
   621 :  data=8'd230   ;
   622 :  data=8'd229   ;
   623 :  data=8'd229   ;
   624 :  data=8'd228   ;
   625 :  data=8'd228   ;
   626 :  data=8'd228   ;
   627 :  data=8'd227   ;
   628 :  data=8'd227   ;
   629 :  data=8'd226   ;
   630 :  data=8'd226   ;
   631 :  data=8'd225   ;
   632 :  data=8'd225   ;
   633 :  data=8'd224   ;
   634 :  data=8'd224   ;
   635 :  data=8'd223   ;
   636 :  data=8'd223   ;
   637 :  data=8'd222   ;
   638 :  data=8'd222   ;
   639 :  data=8'd221   ;
   640 :  data=8'd221   ;
   641 :  data=8'd220   ;
   642 :  data=8'd220   ;
   643 :  data=8'd219   ;
   644 :  data=8'd219   ;
   645 :  data=8'd218   ;
   646 :  data=8'd218   ;
   647 :  data=8'd217   ;
   648 :  data=8'd216   ;
   649 :  data=8'd216   ;
   650 :  data=8'd215   ;
   651 :  data=8'd215   ;
   652 :  data=8'd214   ;
   653 :  data=8'd214   ;
   654 :  data=8'd213   ;
   655 :  data=8'd213   ;
   656 :  data=8'd212   ;
   657 :  data=8'd212   ;
   658 :  data=8'd211   ;
   659 :  data=8'd210   ;
   660 :  data=8'd210   ;
   661 :  data=8'd209   ;
   662 :  data=8'd209   ;
   663 :  data=8'd208   ;
   664 :  data=8'd208   ;
   665 :  data=8'd207   ;
   666 :  data=8'd206   ;
   667 :  data=8'd206   ;
   668 :  data=8'd205   ;
   669 :  data=8'd205   ;
   670 :  data=8'd204   ;
   671 :  data=8'd203   ;
   672 :  data=8'd203   ;
   673 :  data=8'd202   ;
   674 :  data=8'd202   ;
   675 :  data=8'd201   ;
   676 :  data=8'd200   ;
   677 :  data=8'd200   ;
   678 :  data=8'd199   ;
   679 :  data=8'd198   ;
   680 :  data=8'd198   ;
   681 :  data=8'd197   ;
   682 :  data=8'd197   ;
   683 :  data=8'd196   ;
   684 :  data=8'd195   ;
   685 :  data=8'd195   ;
   686 :  data=8'd194   ;
   687 :  data=8'd193   ;
   688 :  data=8'd193   ;
   689 :  data=8'd192   ;
   690 :  data=8'd192   ;
   691 :  data=8'd191   ;
   692 :  data=8'd190   ;
   693 :  data=8'd190   ;
   694 :  data=8'd189   ;
   695 :  data=8'd188   ;
   696 :  data=8'd188   ;
   697 :  data=8'd187   ;
   698 :  data=8'd186   ;
   699 :  data=8'd186   ;
   700 :  data=8'd185   ;
   701 :  data=8'd184   ;
   702 :  data=8'd184   ;
   703 :  data=8'd183   ;
   704 :  data=8'd182   ;
   705 :  data=8'd182   ;
   706 :  data=8'd181   ;
   707 :  data=8'd180   ;
   708 :  data=8'd180   ;
   709 :  data=8'd179   ;
   710 :  data=8'd178   ;
   711 :  data=8'd178   ;
   712 :  data=8'd177   ;
   713 :  data=8'd176   ;
   714 :  data=8'd176   ;
   715 :  data=8'd175   ;
   716 :  data=8'd174   ;
   717 :  data=8'd174   ;
   718 :  data=8'd173   ;
   719 :  data=8'd172   ;
   720 :  data=8'd171   ;
   721 :  data=8'd171   ;
   722 :  data=8'd170   ;
   723 :  data=8'd169   ;
   724 :  data=8'd169   ;
   725 :  data=8'd168   ;
   726 :  data=8'd167   ;
   727 :  data=8'd167   ;
   728 :  data=8'd166   ;
   729 :  data=8'd165   ;
   730 :  data=8'd164   ;
   731 :  data=8'd164   ;
   732 :  data=8'd163   ;
   733 :  data=8'd162   ;
   734 :  data=8'd162   ;
   735 :  data=8'd161   ;
   736 :  data=8'd160   ;
   737 :  data=8'd159   ;
   738 :  data=8'd159   ;
   739 :  data=8'd158   ;
   740 :  data=8'd157   ;
   741 :  data=8'd157   ;
   742 :  data=8'd156   ;
   743 :  data=8'd155   ;
   744 :  data=8'd154   ;
   745 :  data=8'd154   ;
   746 :  data=8'd153   ;
   747 :  data=8'd152   ;
   748 :  data=8'd152   ;
   749 :  data=8'd151   ;
   750 :  data=8'd150   ;
   751 :  data=8'd149   ;
   752 :  data=8'd149   ;
   753 :  data=8'd148   ;
   754 :  data=8'd147   ;
   755 :  data=8'd147   ;
   756 :  data=8'd146   ;
   757 :  data=8'd145   ;
   758 :  data=8'd144   ;
   759 :  data=8'd144   ;
   760 :  data=8'd143   ;
   761 :  data=8'd142   ;
   762 :  data=8'd142   ;
   763 :  data=8'd141   ;
   764 :  data=8'd140   ;
   765 :  data=8'd139   ;
   766 :  data=8'd139   ;
   767 :  data=8'd138   ;
   768 :  data=8'd137   ;
   769 :  data=8'd136   ;
   770 :  data=8'd136   ;
   771 :  data=8'd135   ;
   772 :  data=8'd134   ;
   773 :  data=8'd134   ;
   774 :  data=8'd133   ;
   775 :  data=8'd132   ;
   776 :  data=8'd131   ;
   777 :  data=8'd131   ;
   778 :  data=8'd130   ;
   779 :  data=8'd129   ;
   780 :  data=8'd129   ;
   781 :  data=8'd128   ;
   782 :  data=8'd127   ;
   783 :  data=8'd126   ;
   784 :  data=8'd126   ;
   785 :  data=8'd125   ;
   786 :  data=8'd124   ;
   787 :  data=8'd123   ;
   788 :  data=8'd123   ;
   789 :  data=8'd122   ;
   790 :  data=8'd121   ;
   791 :  data=8'd121   ;
   792 :  data=8'd120   ;
   793 :  data=8'd119   ;
   794 :  data=8'd118   ;
   795 :  data=8'd118   ;
   796 :  data=8'd117   ;
   797 :  data=8'd116   ;
   798 :  data=8'd116   ;
   799 :  data=8'd115   ;
   800 :  data=8'd114   ;
   801 :  data=8'd114   ;
   802 :  data=8'd113   ;
   803 :  data=8'd112   ;
   804 :  data=8'd111   ;
   805 :  data=8'd111   ;
   806 :  data=8'd110   ;
   807 :  data=8'd109   ;
   808 :  data=8'd109   ;
   809 :  data=8'd108   ;
   810 :  data=8'd107   ;
   811 :  data=8'd106   ;
   812 :  data=8'd106   ;
   813 :  data=8'd105   ;
   814 :  data=8'd104   ;
   815 :  data=8'd104   ;
   816 :  data=8'd103   ;
   817 :  data=8'd102   ;
   818 :  data=8'd102   ;
   819 :  data=8'd101   ;
   820 :  data=8'd100   ;
   821 :  data=8'd100   ;
   822 :  data=8'd99    ;
   823 :  data=8'd98    ;
   824 :  data=8'd98    ;
   825 :  data=8'd97    ;
   826 :  data=8'd96    ;
   827 :  data=8'd95    ;
   828 :  data=8'd95    ;
   829 :  data=8'd94    ;
   830 :  data=8'd93    ;
   831 :  data=8'd93    ;
   832 :  data=8'd92    ;
   833 :  data=8'd91    ;
   834 :  data=8'd91    ;
   835 :  data=8'd90    ;
   836 :  data=8'd89    ;
   837 :  data=8'd89    ;
   838 :  data=8'd88    ;
   839 :  data=8'd88    ;
   840 :  data=8'd87    ;
   841 :  data=8'd86    ;
   842 :  data=8'd86    ;
   843 :  data=8'd85    ;
   844 :  data=8'd84    ;
   845 :  data=8'd84    ;
   846 :  data=8'd83    ;
   847 :  data=8'd82    ;
   848 :  data=8'd82    ;
   849 :  data=8'd81    ;
   850 :  data=8'd80    ;
   851 :  data=8'd80    ;
   852 :  data=8'd79    ;
   853 :  data=8'd79    ;
   854 :  data=8'd78    ;
   855 :  data=8'd77    ;
   856 :  data=8'd77    ;
   857 :  data=8'd76    ;
   858 :  data=8'd75    ;
   859 :  data=8'd75    ;
   860 :  data=8'd74    ;
   861 :  data=8'd74    ;
   862 :  data=8'd73    ;
   863 :  data=8'd72    ;
   864 :  data=8'd72    ;
   865 :  data=8'd71    ;
   866 :  data=8'd71    ;
   867 :  data=8'd70    ;
   868 :  data=8'd69    ;
   869 :  data=8'd69    ;
   870 :  data=8'd68    ;
   871 :  data=8'd68    ;
   872 :  data=8'd67    ;
   873 :  data=8'd67    ;
   874 :  data=8'd66    ;
   875 :  data=8'd65    ;
   876 :  data=8'd65    ;
   877 :  data=8'd64    ;
   878 :  data=8'd64    ;
   879 :  data=8'd63    ;
   880 :  data=8'd63    ;
   881 :  data=8'd62    ;
   882 :  data=8'd61    ;
   883 :  data=8'd61    ;
   884 :  data=8'd60    ;
   885 :  data=8'd60    ;
   886 :  data=8'd59    ;
   887 :  data=8'd59    ;
   888 :  data=8'd58    ;
   889 :  data=8'd58    ;
   890 :  data=8'd57    ;
   891 :  data=8'd57    ;
   892 :  data=8'd56    ;
   893 :  data=8'd56    ;
   894 :  data=8'd55    ;
   895 :  data=8'd55    ;
   896 :  data=8'd54    ;
   897 :  data=8'd54    ;
   898 :  data=8'd53    ;
   899 :  data=8'd53    ;
   900 :  data=8'd52    ;
   901 :  data=8'd52    ;
   902 :  data=8'd51    ;
   903 :  data=8'd51    ;
   904 :  data=8'd50    ;
   905 :  data=8'd50    ;
   906 :  data=8'd49    ;
   907 :  data=8'd49    ;
   908 :  data=8'd48    ;
   909 :  data=8'd48    ;
   910 :  data=8'd47    ;
   911 :  data=8'd47    ;
   912 :  data=8'd46    ;
   913 :  data=8'd46    ;
   914 :  data=8'd45    ;
   915 :  data=8'd45    ;
   916 :  data=8'd45    ;
   917 :  data=8'd44    ;
   918 :  data=8'd44    ;
   919 :  data=8'd43    ;
   920 :  data=8'd43    ;
   921 :  data=8'd42    ;
   922 :  data=8'd42    ;
   923 :  data=8'd42    ;
   924 :  data=8'd41    ;
   925 :  data=8'd41    ;
   926 :  data=8'd40    ;
   927 :  data=8'd40    ;
   928 :  data=8'd39    ;
   929 :  data=8'd39    ;
   930 :  data=8'd39    ;
   931 :  data=8'd38    ;
   932 :  data=8'd38    ;
   933 :  data=8'd38    ;
   934 :  data=8'd37    ;
   935 :  data=8'd37    ;
   936 :  data=8'd36    ;
   937 :  data=8'd36    ;
   938 :  data=8'd36    ;
   939 :  data=8'd35    ;
   940 :  data=8'd35    ;
   941 :  data=8'd35    ;
   942 :  data=8'd34    ;
   943 :  data=8'd34    ;
   944 :  data=8'd34    ;
   945 :  data=8'd33    ;
   946 :  data=8'd33    ;
   947 :  data=8'd33    ;
   948 :  data=8'd32    ;
   949 :  data=8'd32    ;
   950 :  data=8'd32    ;
   951 :  data=8'd31    ;
   952 :  data=8'd31    ;
   953 :  data=8'd31    ;
   954 :  data=8'd30    ;
   955 :  data=8'd30    ;
   956 :  data=8'd30    ;
   957 :  data=8'd30    ;
   958 :  data=8'd29    ;
   959 :  data=8'd29    ;
   960 :  data=8'd29    ;
   961 :  data=8'd28    ;
   962 :  data=8'd28    ;
   963 :  data=8'd28    ;
   964 :  data=8'd28    ;
   965 :  data=8'd27    ;
   966 :  data=8'd27    ;
   967 :  data=8'd27    ;
   968 :  data=8'd27    ;
   969 :  data=8'd26    ;
   970 :  data=8'd26    ;
   971 :  data=8'd26    ;
   972 :  data=8'd26    ;
   973 :  data=8'd25    ;
   974 :  data=8'd25    ;
   975 :  data=8'd25    ;
   976 :  data=8'd25    ;
   977 :  data=8'd25    ;
   978 :  data=8'd24    ;
   979 :  data=8'd24    ;
   980 :  data=8'd24    ;
   981 :  data=8'd24    ;
   982 :  data=8'd24    ;
   983 :  data=8'd24    ;
   984 :  data=8'd23    ;
   985 :  data=8'd23    ;
   986 :  data=8'd23    ;
   987 :  data=8'd23    ;
   988 :  data=8'd23    ;
   989 :  data=8'd23    ;
   990 :  data=8'd22    ;
   991 :  data=8'd22    ;
   992 :  data=8'd22    ;
   993 :  data=8'd22    ;
   994 :  data=8'd22    ;
   995 :  data=8'd22    ;
   996 :  data=8'd22    ;
   997 :  data=8'd21    ;
   998 :  data=8'd21    ;
   999 :  data=8'd21    ;
   1000 : data=8'd21    ;
   1001 : data=8'd21    ;
   1002 : data=8'd21    ;
   1003 : data=8'd21    ;
   1004 : data=8'd21    ;
   1005 : data=8'd21    ;
   1006 : data=8'd21    ;
   1007 : data=8'd21    ;
   1008 : data=8'd20    ;
   1009 : data=8'd20    ;
   1010 : data=8'd20    ;
   1011 : data=8'd20    ;
   1012 : data=8'd20    ;
   1013 : data=8'd20    ;
   1014 : data=8'd10    ;
   1015 : data=8'd10    ;
   1016 : data=8'd10    ;
   1017 : data=8'd10    ;
   1018 : data=8'd10    ;
   1019 : data=8'd10    ;
   1020 : data=8'd0    ;
   1021 : data=8'd0    ;
   1022 : data=8'd0    ;
   1023 : data=8'd0    ;
               
      default:                 
            data=    'd0;     

endcase

end






endmodule