module d(
        input wire [10:0]i,
        output reg [31:0] data
   );
always @(*) begin
case(i)
   0 :   data= -1921  ;
   1 :   data= -1932  ;
   2 :   data= -1938  ;
   3 :   data= -1965  ;
   4 :   data= -1985  ;
   5 :   data= -1977  ;
   6 :   data= -2002  ;
   7 :   data= -2051  ;
   8 :   data= -2024  ;
   9 :   data= -1945  ;
   10 :  data= -1932  ;
   11 :  data= -1971  ;
   12 :  data= -1953  ;
   13 :  data= -1893  ;
   14 :  data= -1900  ;
   15 :  data= -1960  ;
   16 :  data= -1954  ;
   17 :  data= -1874  ;
   18 :  data= -1816  ;
   19 :  data= -1803  ;
   20 :  data= -1783  ;
   21 :  data= -1747  ;
   22 :  data= -1712  ;
   23 :  data= -1649  ;
   24 :  data= -1554  ;
   25 :  data= -1501  ;
   26 :  data= -1518  ;
   27 :  data= -1539  ;
   28 :  data= -1533  ;
   29 :  data= -1530  ;
   30 :  data= -1508  ;
   31 :  data= -1448  ;
   32 :  data= -1409  ;
   33 :  data= -1414  ;
   34 :  data= -1415  ;
   35 :  data= -1391  ;
   36 :  data= -1333  ;
   37 :  data= -1243  ;
   38 :  data= -1184  ;
   39 :  data= -1163  ;
   40 :  data= -1111  ;
   41 :  data= -1071  ;
   42 :  data= -1097  ;
   43 :  data= -1068  ;
   44 :  data= -946  ;
   45 :  data= -891  ;
   46 :  data= -917  ;
   47 :  data= -889  ;
   48 :  data= -853  ;
   49 :  data= -922  ;
   50 :  data= -1007  ;
   51 :  data= -990  ;
   52 :  data= -927  ;
   53 :  data= -909  ;
   54 :  data= -929  ;
   55 :  data= -931  ;
   56 :  data= -904  ;
   57 :  data= -911  ;
   58 :  data= -970  ;
   59 :  data= -1001  ;
   60 :  data= -981  ;
   61 :  data= -997  ;
   62 :  data= -1070  ;
   63 :  data= -1103  ;
   64 :  data= -1071  ;
   65 :  data= -1061  ;
   66 :  data= -1109  ;
   67 :  data= -1173  ;
   68 :  data= -1221  ;
   69 :  data= -1265  ;
   70 :  data= -1316  ;
   71 :  data= -1352  ;
   72 :  data= -1356  ;
   73 :  data= -1352  ;
   74 :  data= -1357  ;
   75 :  data= -1329  ;
   76 :  data= -1281  ;
   77 :  data= -1289  ;
   78 :  data= -1320  ;
   79 :  data= -1279  ;
   80 :  data= -1227  ;
   81 :  data= -1255  ;
   82 :  data= -1287  ;
   83 :  data= -1273  ;
   84 :  data= -1286  ;
   85 :  data= -1328  ;
   86 :  data= -1307  ;
   87 :  data= -1235  ;
   88 :  data= -1199  ;
   89 :  data= -1227  ;
   90 :  data= -1265  ;
   91 :  data= -1240  ;
   92 :  data= -1177  ;
   93 :  data= -1165  ;
   94 :  data= -1203  ;
   95 :  data= -1209  ;
   96 :  data= -1188  ;
   97 :  data= -1172  ;
   98 :  data= -1138  ;
   99 :  data= -1096  ;
   100 :  data=-1094  ;
   101 :  data=-1115  ;
   102 :  data=-1122  ;
   103 :  data=-1119  ;
   104 :  data=-1101  ;
   105 :  data=-1063  ;
   106 :  data=-1025  ;
   107 :  data=-972  ;
   108 :  data=-890  ;
   109 :  data=-815  ;
   110 :  data=-781  ;
   111 :  data=-779  ;
   112 :  data=-789  ;
   113 :  data=-783  ;
   114 :  data=-750  ;
   115 :  data=-748  ;
   116 :  data=-778  ;
   117 :  data=-741  ;
   118 :  data=-665  ;
   119 :  data=-691  ;
   120 :  data=-771  ;
   121 :  data=-748  ;
   122 :  data=-665  ;
   123 :  data=-644  ;
   124 :  data=-637  ;
   125 :  data=-590  ;
   126 :  data=-563  ;
   127 :  data=-565  ;
   128 :  data=-543  ;
   129 :  data=-511  ;
   130 :  data=-515  ;
   131 :  data=-542  ;
   132 :  data=-536  ;
   133 :  data=-472  ;
   134 :  data=-426  ;
   135 :  data=-481  ;
   136 :  data=-545  ;
   137 :  data=-493  ;
   138 :  data=-410  ;
   139 :  data=-395  ;
   140 :  data=-356  ;
   141 :  data=-239  ;
   142 :  data=-161  ;
   143 :  data=-149  ;
   144 :  data=-102  ;
   145 :  data=-3  ;
   146 :  data=79  ;
   147 :  data=118  ;
   148 :  data=133  ;
   149 :  data=179  ;
   150 :  data=258  ;
   151 :  data=285  ;
   152 :  data=243  ;
   153 :  data=243  ;
   154 :  data=302  ;
   155 :  data=318  ;
   156 :  data=290  ;
   157 :  data=292  ;
   158 :  data=310  ;
   159 :  data=308  ;
   160 :  data=312  ;
   161 :  data=327  ;
   162 :  data=332  ;
   163 :  data=315  ;
   164 :  data=281  ;
   165 :  data=257  ;
   166 :  data=271  ;
   167 :  data=297  ;
   168 :  data=290  ;
   169 :  data=253  ;
   170 :  data=195  ;
   171 :  data=150  ;
   172 :  data=174  ;
   173 :  data=235  ;
   174 :  data=239  ;
   175 :  data=199  ;
   176 :  data=193  ;
   177 :  data=217  ;
   178 :  data=220  ;
   179 :  data=199  ;
   180 :  data=175  ;
   181 :  data=161  ;
   182 :  data=150  ;
   183 :  data=129  ;
   184 :  data=111  ;
   185 :  data=113  ;
   186 :  data=110  ;
   187 :  data=117  ;
   188 :  data=185  ;
   189 :  data=255  ;
   190 :  data=233  ;
   191 :  data=195  ;
   192 :  data=230  ;
   193 :  data=246  ;
   194 :  data=190  ;
   195 :  data=178  ;
   196 :  data=240  ;
   197 :  data=267  ;
   198 :  data=228  ;
   199 :  data=180  ;
   200 :  data=149  ;
   201 :  data=131  ;
   202 :  data=105  ;
   203 :  data=49  ;
   204 :  data=1  ;
   205 :  data=-9  ;
   206 :  data=-6  ;
   207 :  data=31  ;
   208 :  data=118  ;
   209 :  data=151  ;
   210 :  data=112  ;
   211 :  data=137  ;
   212 :  data=227  ;
   213 :  data=257  ;
   214 :  data=265  ;
   215 :  data=355  ;
   216 :  data=441  ;
   217 :  data=438  ;
   218 :  data=438  ;
   219 :  data=506  ;
   220 :  data=557  ;
   221 :  data=531  ;
   222 :  data=507  ;
   223 :  data=568  ;
   224 :  data=679  ;
   225 :  data=740  ;
   226 :  data=736  ;
   227 :  data=741  ;
   228 :  data=797  ;
   229 :  data=863  ;
   230 :  data=899  ;
   231 :  data=906  ;
   232 :  data=909  ;
   233 :  data=930  ;
   234 :  data=962  ;
   235 :  data=974  ;
   236 :  data=952  ;
   237 :  data=917  ;
   238 :  data=884  ;
   239 :  data=853  ;
   240 :  data=846  ;
   241 :  data=855  ;
   242 :  data=828  ;
   243 :  data=771  ;
   244 :  data=747  ;
   245 :  data=742  ;
   246 :  data=699  ;
   247 :  data=632  ;
   248 :  data=580  ;
   249 :  data=541  ;
   250 :  data=509  ;
   251 :  data=476  ;
   252 :  data=436  ;
   253 :  data=422  ;
   254 :  data=445  ;
   255 :  data=451  ;
   256 :  data=409  ;
   257 :  data=362  ;
   258 :  data=352  ;
   259 :  data=354  ;
   260 :  data=322  ;
   261 :  data=266  ;
   262 :  data=229  ;
   263 :  data=206  ;
   264 :  data=157  ;
   265 :  data=92  ;
   266 :  data=26  ;
   267 :  data=-35  ;
   268 :  data=-63  ;
   269 :  data=-50  ;
   270 :  data=-60  ;
   271 :  data=-96  ;
   272 :  data=-93  ;
   273 :  data=-62  ;
   274 :  data=-55  ;
   275 :  data=-56  ;
   276 :  data=-45  ;
   277 :  data=-25  ;
   278 :  data=31  ;
   279 :  data=115  ;
   280 :  data=159  ;
   281 :  data=165  ;
   282 :  data=197  ;
   283 :  data=241  ;
   284 :  data=243  ;
   285 :  data=242  ;
   286 :  data=296  ;
   287 :  data=339  ;
   288 :  data=305  ;
   289 :  data=282  ;
   290 :  data=341  ;
   291 :  data=379  ;
   292 :  data=326  ;
   293 :  data=301  ;
   294 :  data=370  ;
   295 :  data=425  ;
   296 :  data=416  ;
   297 :  data=444  ;
   298 :  data=539  ;
   299 :  data=588  ;
   300 :  data=548  ;
   301 :  data=531  ;
   302 :  data=607  ;
   303 :  data=706  ;
   304 :  data=761  ;
   305 :  data=797  ;
   306 :  data=830  ;
   307 :  data=817  ;
   308 :  data=772  ;
   309 :  data=772  ;
   310 :  data=817  ;
   311 :  data=829  ;
   312 :  data=821  ;
   313 :  data=867  ;
   314 :  data=918  ;
   315 :  data=900  ;
   316 :  data=892  ;
   317 :  data=972  ;
   318 :  data=1044  ;
   319 :  data=1045  ;
   320 :  data=1064  ;
   321 :  data=1129  ;
   322 :  data=1153  ;
   323 :  data=1128  ;
   324 :  data=1127  ;
   325 :  data=1157  ;
   326 :  data=1158  ;
   327 :  data=1101  ;
   328 :  data=1029  ;
   329 :  data=972  ;
   330 :  data=903  ;
   331 :  data=830  ;
   332 :  data=807  ;
   333 :  data=794  ;
   334 :  data=723  ;
   335 :  data=648  ;
   336 :  data=628  ;
   337 :  data=601  ;
   338 :  data=542  ;
   339 :  data=512  ;
   340 :  data=516  ;
   341 :  data=492  ;
   342 :  data=429  ;
   343 :  data=374  ;
   344 :  data=364  ;
   345 :  data=378  ;
   346 :  data=361  ;
   347 :  data=325  ;
   348 :  data=319  ;
   349 :  data=320  ;
   350 :  data=302  ;
   351 :  data=289  ;
   352 :  data=272  ;
   353 :  data=218  ;
   354 :  data=178  ;
   355 :  data=210  ;
   356 :  data=252  ;
   357 :  data=249  ;
   358 :  data=255  ;
   359 :  data=285  ;
   360 :  data=282  ;
   361 :  data=269  ;
   362 :  data=307  ;
   363 :  data=343  ;
   364 :  data=330  ;
   365 :  data=332  ;
   366 :  data=363  ;
   367 :  data=350  ;
   368 :  data=326  ;
   369 :  data=380  ;
   370 :  data=462  ;
   371 :  data=457  ;
   372 :  data=386  ;
   373 :  data=353  ;
   374 :  data=380  ;
   375 :  data=395  ;
   376 :  data=373  ;
   377 :  data=355  ;
   378 :  data=342  ;
   379 :  data=302  ;
   380 :  data=271  ;
   381 :  data=289  ;
   382 :  data=323  ;
   383 :  data=357  ;
   384 :  data=404  ;
   385 :  data=421  ;
   386 :  data=391  ;
   387 :  data=390  ;
   388 :  data=451  ;
   389 :  data=507  ;
   390 :  data=526  ;
   391 :  data=540  ;
   392 :  data=546  ;
   393 :  data=501  ;
   394 :  data=404  ;
   395 :  data=339  ;
   396 :  data=370  ;
   397 :  data=426  ;
   398 :  data=413  ;
   399 :  data=373  ;
   400 :  data=385  ;
   401 :  data=399  ;
   402 :  data=366  ;
   403 :  data=357  ;
   404 :  data=405  ;
   405 :  data=426  ;
   406 :  data=392  ;
   407 :  data=360  ;
   408 :  data=317  ;
   409 :  data=237  ;
   410 :  data=202  ;
   411 :  data=256  ;
   412 :  data=292  ;
   413 :  data=249  ;
   414 :  data=228  ;
   415 :  data=292  ;
   416 :  data=355  ;
   417 :  data=354  ;
   418 :  data=364  ;
   419 :  data=443  ;
   420 :  data=504  ;
   421 :  data=504  ;
   422 :  data=533  ;
   423 :  data=607  ;
   424 :  data=633  ;
   425 :  data=643  ;
   426 :  data=712  ;
   427 :  data=749  ;
   428 :  data=708  ;
   429 :  data=724  ;
   430 :  data=825  ;
   431 :  data=870  ;
   432 :  data=842  ;
   433 :  data=842  ;
   434 :  data=878  ;
   435 :  data=901  ;
   436 :  data=905  ;
   437 :  data=904  ;
   438 :  data=932  ;
   439 :  data=1002  ;
   440 :  data=1052  ;
   441 :  data=1028  ;
   442 :  data=974  ;
   443 :  data=957  ;
   444 :  data=974  ;
   445 :  data=990  ;
   446 :  data=997  ;
   447 :  data=1011  ;
   448 :  data=1034  ;
   449 :  data=1018  ;
   450 :  data=942  ;
   451 :  data=872  ;
   452 :  data=885  ;
   453 :  data=955  ;
   454 :  data=1002  ;
   455 :  data=1019  ;
   456 :  data=1050  ;
   457 :  data=1093  ;
   458 :  data=1098  ;
   459 :  data=1059  ;
   460 :  data=1025  ;
   461 :  data=1023  ;
   462 :  data=1024  ;
   463 :  data=1005  ;
   464 :  data=972  ;
   465 :  data=941  ;
   466 :  data=927  ;
   467 :  data=934  ;
   468 :  data=932  ;
   469 :  data=905  ;
   470 :  data=877  ;
   471 :  data=855  ;
   472 :  data=823  ;
   473 :  data=789  ;
   474 :  data=762  ;
   475 :  data=719  ;
   476 :  data=679  ;
   477 :  data=675  ;
   478 :  data=655  ;
   479 :  data=585  ;
   480 :  data=549  ;
   481 :  data=584  ;
   482 :  data=611  ;
   483 :  data=611  ;
   484 :  data=639  ;
   485 :  data=695  ;
   486 :  data=757  ;
   487 :  data=814  ;
   488 :  data=830  ;
   489 :  data=822  ;
   490 :  data=879  ;
   491 :  data=980  ;
   492 :  data=1023  ;
   493 :  data=1047  ;
   494 :  data=1122  ;
   495 :  data=1148  ;
   496 :  data=1069  ;
   497 :  data=1036  ;
   498 :  data=1120  ;
   499 :  data=1198  ;
   500 :  data=1238  ;
   501 :  data=1332  ;
   502 :  data=1439  ;
   503 :  data=1451  ;
   504 :  data=1413  ;
   505 :  data=1430  ;
   506 :  data=1483  ;
   507 :  data=1497  ;
   508 :  data=1488  ;
   509 :  data=1515  ;
   510 :  data=1563  ;
   511 :  data=1575  ;
   512 :  data=1566  ;
   513 :  data=1584  ;
   514 :  data=1597  ;
   515 :  data=1558  ;
   516 :  data=1510  ;
   517 :  data=1510  ;
   518 :  data=1539  ;
   519 :  data=1564  ;
   520 :  data=1586  ;
   521 :  data=1595  ;
   522 :  data=1584  ;
   523 :  data=1563  ;
   524 :  data=1540  ;
   525 :  data=1526  ;
   526 :  data=1519  ;
   527 :  data=1497  ;
   528 :  data=1463  ;
   529 :  data=1439  ;
   530 :  data=1397  ;
   531 :  data=1320  ;
   532 :  data=1257  ;
   533 :  data=1235  ;
   534 :  data=1209  ;
   535 :  data=1158  ;
   536 :  data=1087  ;
   537 :  data=982  ;
   538 :  data=873  ;
   539 :  data=824  ;
   540 :  data=809  ;
   541 :  data=767  ;
   542 :  data=708  ;
   543 :  data=650  ;
   544 :  data=573  ;
   545 :  data=515  ;
   546 :  data=515  ;
   547 :  data=517  ;
   548 :  data=482  ;
   549 :  data=463  ;
   550 :  data=485  ;
   551 :  data=492  ;
   552 :  data=463  ;
   553 :  data=433  ;
   554 :  data=420  ;
   555 :  data=419  ;
   556 :  data=425  ;
   557 :  data=437  ;
   558 :  data=464  ;
   559 :  data=501  ;
   560 :  data=501  ;
   561 :  data=455  ;
   562 :  data=431  ;
   563 :  data=470  ;
   564 :  data=523  ;
   565 :  data=539  ;
   566 :  data=534  ;
   567 :  data=522  ;
   568 :  data=499  ;
   569 :  data=483  ;
   570 :  data=487  ;
   571 :  data=490  ;
   572 :  data=493  ;
   573 :  data=524  ;
   574 :  data=572  ;
   575 :  data=602  ;
   576 :  data=623  ;
   577 :  data=664  ;
   578 :  data=697  ;
   579 :  data=696  ;
   580 :  data=705  ;
   581 :  data=764  ;
   582 :  data=825  ;
   583 :  data=831  ;
   584 :  data=825  ;
   585 :  data=824  ;
   586 :  data=761  ;
   587 :  data=673  ;
   588 :  data=670  ;
   589 :  data=695  ;
   590 :  data=650  ;
   591 :  data=628  ;
   592 :  data=690  ;
   593 :  data=716  ;
   594 :  data=687  ;
   595 :  data=703  ;
   596 :  data=726  ;
   597 :  data=699  ;
   598 :  data=702  ;
   599 :  data=750  ;
   600 :  data=747  ;
   601 :  data=689  ;
   602 :  data=625  ;
   603 :  data=558  ;
   604 :  data=492  ;
   605 :  data=432  ;
   606 :  data=374  ;
   607 :  data=362  ;
   608 :  data=386  ;
   609 :  data=353  ;
   610 :  data=281  ;
   611 :  data=261  ;
   612 :  data=246  ;
   613 :  data=191  ;
   614 :  data=182  ;
   615 :  data=223  ;
   616 :  data=202  ;
   617 :  data=134  ;
   618 :  data=110  ;
   619 :  data=111  ;
   620 :  data=82  ;
   621 :  data=26  ;
   622 :  data=-33  ;
   623 :  data=-63  ;
   624 :  data=-66  ;
   625 :  data=-72  ;
   626 :  data=-52  ;
   627 :  data=11  ;
   628 :  data=41  ;
   629 :  data=41  ;
   630 :  data=117  ;
   631 :  data=216  ;
   632 :  data=202  ;
   633 :  data=150  ;
   634 :  data=175  ;
   635 :  data=199  ;
   636 :  data=156  ;
   637 :  data=108  ;
   638 :  data=74  ;
   639 :  data=23  ;
   640 :  data=-19  ;
   641 :  data=-18  ;
   642 :  data=34  ;
   643 :  data=138  ;
   644 :  data=225  ;
   645 :  data=237  ;
   646 :  data=236  ;
   647 :  data=282  ;
   648 :  data=325  ;
   649 :  data=308  ;
   650 :  data=239  ;
   651 :  data=129  ;
   652 :  data=-4  ;
   653 :  data=-127  ;
   654 :  data=-218  ;
   655 :  data=-272  ;
   656 :  data=-285  ;
   657 :  data=-288  ;
   658 :  data=-308  ;
   659 :  data=-325  ;
   660 :  data=-305  ;
   661 :  data=-248  ;
   662 :  data=-193  ;
   663 :  data=-193  ;
   664 :  data=-241  ;
   665 :  data=-274  ;
   666 :  data=-294  ;
   667 :  data=-379  ;
   668 :  data=-531  ;
   669 :  data=-657  ;
   670 :  data=-720  ;
   671 :  data=-742  ;
   672 :  data=-724  ;
   673 :  data=-696  ;
   674 :  data=-702  ;
   675 :  data=-719  ;
   676 :  data=-727  ;
   677 :  data=-762  ;
   678 :  data=-788  ;
   679 :  data=-744  ;
   680 :  data=-714  ;
   681 :  data=-774  ;
   682 :  data=-830  ;
   683 :  data=-823  ;
   684 :  data=-821  ;
   685 :  data=-829  ;
   686 :  data=-813  ;
   687 :  data=-827  ;
   688 :  data=-869  ;
   689 :  data=-835  ;
   690 :  data=-740  ;
   691 :  data=-693  ;
   692 :  data=-671  ;
   693 :  data=-605  ;
   694 :  data=-521  ;
   695 :  data=-444  ;
   696 :  data=-355  ;
   697 :  data=-274  ;
   698 :  data=-214  ;
   699 :  data=-141  ;
   700 :  data=-49  ;
   701 :  data=19  ;
   702 :  data=55  ;
   703 :  data=66  ;
   704 :  data=56  ;
   705 :  data=47  ;
   706 :  data=34  ;
   707 :  data=-17  ;
   708 :  data=-63  ;
   709 :  data=-18  ;
   710 :  data=72  ;
   711 :  data=118  ;
   712 :  data=175  ;
   713 :  data=296  ;
   714 :  data=358  ;
   715 :  data=296  ;
   716 :  data=255  ;
   717 :  data=314  ;
   718 :  data=352  ;
   719 :  data=323  ;
   720 :  data=325  ;
   721 :  data=351  ;
   722 :  data=285  ;
   723 :  data=139  ;
   724 :  data=40  ;
   725 :  data=15  ;
   726 :  data=14  ;
   727 :  data=49  ;
   728 :  data=123  ;
   729 :  data=151  ;
   730 :  data=101  ;
   731 :  data=48  ;
   732 :  data=20  ;
   733 :  data=-17  ;
   734 :  data=-29  ;
   735 :  data=4  ;
   736 :  data=1  ;
   737 :  data=-61  ;
   738 :  data=-109  ;
   739 :  data=-156  ;
   740 :  data=-253  ;
   741 :  data=-343  ;
   742 :  data=-404  ;
   743 :  data=-495  ;
   744 :  data=-574  ;
   745 :  data=-590  ;
   746 :  data=-637  ;
   747 :  data=-752  ;
   748 :  data=-829  ;
   749 :  data=-855  ;
   750 :  data=-874  ;
   751 :  data=-836  ;
   752 :  data=-786  ;
   753 :  data=-852  ;
   754 :  data=-963  ;
   755 :  data=-983  ;
   756 :  data=-964  ;
   757 :  data=-964  ;
   758 :  data=-955  ;
   759 :  data=-989  ;
   760 :  data=-1087  ;
   761 :  data=-1123  ;
   762 :  data=-1051  ;
   763 :  data=-955  ;
   764 :  data=-871  ;
   765 :  data=-816  ;
   766 :  data=-822  ;
   767 :  data=-819  ;
   768 :  data=-741  ;
   769 :  data=-654  ;
   770 :  data=-618  ;
   771 :  data=-605  ;
   772 :  data=-597  ;
   773 :  data=-588  ;
   774 :  data=-550  ;
   775 :  data=-485  ;
   776 :  data=-397  ;
   777 :  data=-274  ;
   778 :  data=-138  ;
   779 :  data=-30  ;
   780 :  data=45  ;
   781 :  data=101  ;
   782 :  data=157  ;
   783 :  data=231  ;
   784 :  data=275  ;
   785 :  data=255  ;
   786 :  data=227  ;
   787 :  data=215  ;
   788 :  data=186  ;
   789 :  data=181  ;
   790 :  data=231  ;
   791 :  data=273  ;
   792 :  data=303  ;
   793 :  data=370  ;
   794 :  data=401  ;
   795 :  data=346  ;
   796 :  data=342  ;
   797 :  data=440  ;
   798 :  data=476  ;
   799 :  data=402  ;
   800 :  data=356  ;
   801 :  data=383  ;
   802 :  data=410  ;
   803 :  data=440  ;
   804 :  data=515  ;
   805 :  data=587  ;
   806 :  data=587  ;
   807 :  data=503  ;
   808 :  data=362  ;
   809 :  data=215  ;
   810 :  data=146  ;
   811 :  data=194  ;
   812 :  data=272  ;
   813 :  data=258  ;
   814 :  data=177  ;
   815 :  data=142  ;
   816 :  data=132  ;
   817 :  data=41  ;
   818 :  data=-78  ;
   819 :  data=-91  ;
   820 :  data=-43  ;
   821 :  data=-68  ;
   822 :  data=-151  ;
   823 :  data=-218  ;
   824 :  data=-290  ;
   825 :  data=-386  ;
   826 :  data=-454  ;
   827 :  data=-480  ;
   828 :  data=-457  ;
   829 :  data=-351  ;
   830 :  data=-223  ;
   831 :  data=-173  ;
   832 :  data=-156  ;
   833 :  data=-103  ;
   834 :  data=-68  ;
   835 :  data=-70  ;
   836 :  data=-33  ;
   837 :  data=23  ;
   838 :  data=20  ;
   839 :  data=-14  ;
   840 :  data=-19  ;
   841 :  data=0  ;
   842 :  data=41  ;
   843 :  data=110  ;
   844 :  data=175  ;
   845 :  data=226  ;
   846 :  data=285  ;
   847 :  data=336  ;
   848 :  data=353  ;
   849 :  data=330  ;
   850 :  data=268  ;
   851 :  data=228  ;
   852 :  data=274  ;
   853 :  data=356  ;
   854 :  data=409  ;
   855 :  data=473  ;
   856 :  data=562  ;
   857 :  data=610  ;
   858 :  data=637  ;
   859 :  data=706  ;
   860 :  data=754  ;
   861 :  data=719  ;
   862 :  data=688  ;
   863 :  data=714  ;
   864 :  data=718  ;
   865 :  data=674  ;
   866 :  data=669  ;
   867 :  data=726  ;
   868 :  data=789  ;
   869 :  data=833  ;
   870 :  data=867  ;
   871 :  data=882  ;
   872 :  data=856  ;
   873 :  data=803  ;
   874 :  data=784  ;
   875 :  data=833  ;
   876 :  data=888  ;
   877 :  data=864  ;
   878 :  data=794  ;
   879 :  data=766  ;
   880 :  data=771  ;
   881 :  data=741  ;
   882 :  data=698  ;
   883 :  data=708  ;
   884 :  data=736  ;
   885 :  data=705  ;
   886 :  data=639  ;
   887 :  data=592  ;
   888 :  data=523  ;
   889 :  data=377  ;
   890 :  data=230  ;
   891 :  data=156  ;
   892 :  data=85  ;
   893 :  data=-25  ;
   894 :  data=-66  ;
   895 :  data=-1  ;
   896 :  data=13  ;
   897 :  data=-77  ;
   898 :  data=-123  ;
   899 :  data=-70  ;
   900 :  data=-42  ;
   901 :  data=-74  ;
   902 :  data=-83  ;
   903 :  data=-90  ;
   904 :  data=-174  ;
   905 :  data=-321  ;
   906 :  data=-457  ;
   907 :  data=-548  ;
   908 :  data=-594  ;
   909 :  data=-601  ;
   910 :  data=-582  ;
   911 :  data=-575  ;
   912 :  data=-617  ;
   913 :  data=-665  ;
   914 :  data=-648  ;
   915 :  data=-588  ;
   916 :  data=-560  ;
   917 :  data=-557  ;
   918 :  data=-546  ;
   919 :  data=-540  ;
   920 :  data=-547  ;
   921 :  data=-554  ;
   922 :  data=-561  ;
   923 :  data=-550  ;
   924 :  data=-523  ;
   925 :  data=-547  ;
   926 :  data=-649  ;
   927 :  data=-764  ;
   928 :  data=-837  ;
   929 :  data=-873  ;
   930 :  data=-878  ;
   931 :  data=-877  ;
   932 :  data=-902  ;
   933 :  data=-924  ;
   934 :  data=-902  ;
   935 :  data=-861  ;
   936 :  data=-848  ;
   937 :  data=-852  ;
   938 :  data=-834  ;
   939 :  data=-801  ;
   940 :  data=-805  ;
   941 :  data=-860  ;
   942 :  data=-908  ;
   943 :  data=-915  ;
   944 :  data=-932  ;
   945 :  data=-983  ;
   946 :  data=-1020  ;
   947 :  data=-1028  ;
   948 :  data=-1048  ;
   949 :  data=-1080  ;
   950 :  data=-1115  ;
   951 :  data=-1188  ;
   952 :  data=-1284  ;
   953 :  data=-1330  ;
   954 :  data=-1343  ;
   955 :  data=-1407  ;
   956 :  data=-1496  ;
   957 :  data=-1523  ;
   958 :  data=-1516  ;
   959 :  data=-1551  ;
   960 :  data=-1598  ;
   961 :  data=-1594  ;
   962 :  data=-1576  ;
   963 :  data=-1590  ;
   964 :  data=-1598  ;
   965 :  data=-1577  ;
   966 :  data=-1575  ;
   967 :  data=-1629  ;
   968 :  data=-1705  ;
   969 :  data=-1758  ;
   970 :  data=-1780  ;
   971 :  data=-1798  ;
   972 :  data=-1811  ;
   973 :  data=-1789  ;
   974 :  data=-1756  ;
   975 :  data=-1766  ;
   976 :  data=-1791  ;
   977 :  data=-1790  ;
   978 :  data=-1817  ;
   979 :  data=-1888  ;
   980 :  data=-1911  ;
   981 :  data=-1892  ;
   982 :  data=-1941  ;
   983 :  data=-2044  ;
   984 :  data=-2108  ;
   985 :  data=-2141  ;
   986 :  data=-2178  ;
   987 :  data=-2192  ;
   988 :  data=-2176  ;
   989 :  data=-2169  ;
   990 :  data=-2198  ;
   991 :  data=-2264  ;
   992 :  data=-2345  ;
   993 :  data=-2401  ;
   994 :  data=-2435  ;
   995 :  data=-2483  ;
   996 :  data=-2546  ;
   997 :  data=-2591  ;
   998 :  data=-2599  ;
   999 :  data=-2596  ;
   1000 : data=-2607  ;
   1001 : data=-2599  ;
   1002 : data=-2558  ;
   1003 : data=-2564  ;
   1004 : data=-2639  ;
   1005 : data=-2672  ;
   1006 : data=-2623  ;
   1007 : data=-2596  ;
   1008 : data=-2620  ;
   1009 : data=-2643  ;
   1010 : data=-2681  ;
   1011 : data=-2755  ;
   1012 : data=-2809  ;
   1013 : data=-2825  ;
   1014 : data=-2834  ;
   1015 : data=-2819  ;
   1016 : data=-2789  ;
   1017 : data=-2816  ;
   1018 : data=-2904  ;
   1019 : data=-2979  ;
   1020 : data=-3023  ;
   1021 : data=-3070  ;
   1022 : data=-3127  ;
   1023 : data=-3178  ;
   1024 : data=-3209  ;
   1025 : data=-3216  ;
   1026 : data=-3214  ;
   1027 : data=-3221  ;
   1028 : data=-3242  ;
   1029 : data=-3280  ;
   1030 : data=-3320  ;
   1031 : data=-3346  ;
   1032 : data=-3377  ;
   1033 : data=-3421  ;
   1034 : data=-3433  ;
   1035 : data=-3414  ;
   1036 : data=-3420  ;
   1037 : data=-3450  ;
   1038 : data=-3459  ;
   1039 : data=-3451  ;
   1040 : data=-3439  ;
   1041 : data=-3397  ;
   1042 : data=-3337  ;
   1043 : data=-3291  ;
   1044 : data=-3250  ;
   1045 : data=-3197  ;
   1046 : data=-3168  ;
   1047 : data=-3179  ;
   1048 : data=-3193  ;
   1049 : data=-3175  ;
   1050 : data=-3135  ;
   1051 : data=-3102  ;
   1052 : data=-3073  ;
   1053 : data=-3032  ;
   1054 : data=-2995  ;
   1055 : data=-2977  ;
   1056 : data=-2972  ;
   1057 : data=-2991  ;
   1058 : data=-3037  ;
   1059 : data=-3051  ;
   1060 : data=-3017  ;
   1061 : data=-3040  ;
   1062 : data=-3155  ;
   1063 : data=-3259  ;
   1064 : data=-3306  ;
   1065 : data=-3342  ;
   1066 : data=-3359  ;
   1067 : data=-3339  ;
   1068 : data=-3327  ;
   1069 : data=-3332  ;
   1070 : data=-3327  ;
   1071 : data=-3345  ;
   1072 : data=-3391  ;
   1073 : data=-3409  ;
   1074 : data=-3416  ;
   1075 : data=-3472  ;
   1076 : data=-3538  ;
   1077 : data=-3557  ;
   1078 : data=-3555  ;
   1079 : data=-3554  ;
   1080 : data=-3547  ;
   1081 : data=-3546  ;
   1082 : data=-3542  ;
   1083 : data=-3520  ;
   1084 : data=-3532  ;
   1085 : data=-3604  ;
   1086 : data=-3671  ;
   1087 : data=-3700  ;
   1088 : data=-3727  ;
   1089 : data=-3754  ;
   1090 : data=-3748  ;
   1091 : data=-3697  ;
   1092 : data=-3628  ;
   1093 : data=-3614  ;
   1094 : data=-3688  ;
   1095 : data=-3767  ;
   1096 : data=-3778  ;
   1097 : data=-3749  ;
   1098 : data=-3716  ;
   1099 : data=-3687  ;
   1100 : data=-3683  ;
   1101 : data=-3681  ;
   1102 : data=-3639  ;
   1103 : data=-3599  ;
   1104 : data=-3596  ;
   1105 : data=-3573  ;
   1106 : data=-3503  ;
   1107 : data=-3431  ;
   1108 : data=-3367  ;
   1109 : data=-3296  ;
   1110 : data=-3215  ;
   1111 : data=-3116  ;
   1112 : data=-3022  ;
   1113 : data=-2980  ;
   1114 : data=-2963  ;
   1115 : data=-2933  ;
   1116 : data=-2900  ;
   1117 : data=-2843  ;
   1118 : data=-2738  ;
   1119 : data=-2653  ;
   1120 : data=-2611  ;
   1121 : data=-2553  ;
   1122 : data=-2495  ;
   1123 : data=-2481  ;
   1124 : data=-2435  ;
   1125 : data=-2310  ;
   1126 : data=-2175  ;
   1127 : data=-2068  ;
   1128 : data=-1997  ;
   1129 : data=-1997  ;
   1130 : data=-2035  ;
   1131 : data=-2041  ;
   1132 : data=-2023  ;
   1133 : data=-1999  ;
   1134 : data=-1959  ;
   1135 : data=-1929  ;
   1136 : data=-1907  ;
   1137 : data=-1854  ;
   1138 : data=-1816  ;
   1139 : data=-1844  ;
   1140 : data=-1867  ;
   1141 : data=-1839  ;
   1142 : data=-1809  ;
   1143 : data=-1759  ;
   1144 : data=-1648  ;
   1145 : data=-1558  ;
   1146 : data=-1534  ;
   1147 : data=-1504  ;
   1148 : data=-1474  ;
   1149 : data=-1508  ;
   1150 : data=-1538  ;
   1151 : data=-1478  ;
   1152 : data=-1405  ;
   1153 : data=-1401  ;
   1154 : data=-1407  ;
   1155 : data=-1364  ;
   1156 : data=-1307  ;
   1157 : data=-1274  ;
   1158 : data=-1273  ;
   1159 : data=-1324  ;
   1160 : data=-1407  ;
   1161 : data=-1435  ;
   1162 : data=-1366  ;
   1163 : data=-1276  ;
   1164 : data=-1245  ;
   1165 : data=-1241  ;
   1166 : data=-1202  ;
   1167 : data=-1158  ;
   1168 : data=-1183  ;
   1169 : data=-1248  ;
   1170 : data=-1233  ;
   1171 : data=-1097  ;
   1172 : data=-953  ;
   1173 : data=-903  ;
   1174 : data=-912  ;
   1175 : data=-897  ;
   1176 : data=-835  ;
   1177 : data=-767  ;
   1178 : data=-745  ;
   1179 : data=-737  ;
   1180 : data=-639  ;
   1181 : data=-469  ;
   1182 : data=-400  ;
   1183 : data=-461  ;
   1184 : data=-456  ;
   1185 : data=-318  ;
   1186 : data=-202  ;
   1187 : data=-158  ;
   1188 : data=-75  ;
   1189 : data=73  ;
   1190 : data=217  ;
   1191 : data=328  ;
   1192 : data=386  ;
   1193 : data=375  ;
   1194 : data=386  ;
   1195 : data=499  ;
   1196 : data=620  ;
   1197 : data=637  ;
   1198 : data=609  ;
   1199 : data=637  ;
               
      default:                 
            data=    'd0;     

endcase

end



endmodule


